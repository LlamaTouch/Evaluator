[
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      1
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "android:id/parentPanel",
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/customPanel",
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      6
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": "android:id/custom",
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        569
      ],
      [
        922,
        1286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      7
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "765*717",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        584
      ],
      [
        907,
        1271
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*687",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        584
      ],
      [
        907,
        1271
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      9,
      12,
      16
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 7,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*687",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        584
      ],
      [
        907,
        737
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*153",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        584
      ],
      [
        907,
        737
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 9,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*153",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        636
      ],
      [
        694,
        706
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 10,
    "resource_id": "com.google.android.apps.maps:id/dialog_title",
    "scrollable": false,
    "selected": false,
    "size": "470*70",
    "temp_id": 11,
    "text": "Timeline data deleted",
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        737
      ],
      [
        907,
        957
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      13
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*220",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        737
      ],
      [
        907,
        957
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 12,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*220",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        737
      ],
      [
        907,
        957
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*220",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        737
      ],
      [
        855,
        957
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": "com.google.android.apps.maps:id/dialog_body_text",
    "scrollable": false,
    "selected": false,
    "size": "631*220",
    "temp_id": 15,
    "text": "You may also want to check your past searches and the content you've browsed in your Timeline and other apps.",
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        957
      ],
      [
        907,
        1271
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      17
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*314",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        988
      ],
      [
        855,
        1240
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "631*252",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        988
      ],
      [
        855,
        1240
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      19,
      21
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "631*252",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        988
      ],
      [
        855,
        1114
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      20
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Done",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/dialog_positive_button",
    "scrollable": false,
    "selected": false,
    "size": "631*126",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        998
      ],
      [
        855,
        1103
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Done",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "631*105",
    "temp_id": 20,
    "text": "Done",
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        1114
      ],
      [
        855,
        1240
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Go to Web & App Activity",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/dialog_negative_button",
    "scrollable": false,
    "selected": false,
    "size": "631*126",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        224,
        1124
      ],
      [
        855,
        1229
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Go to Web & App Activity",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "631*105",
    "temp_id": 22,
    "text": "Go to Web & App Activity",
    "visible": true
  }
]
