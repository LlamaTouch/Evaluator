[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      99
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 2,
    "resource_id": "com.google.android.apps.magazines:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      6
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 4,
    "resource_id": "com.google.android.apps.magazines:id/main_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      7,
      9,
      13
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 5,
    "resource_id": "com.google.android.apps.magazines:id/search_fragment",
    "scrollable": true,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 6,
    "resource_id": "com.google.android.apps.magazines:id/search_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 7,
    "resource_id": "com.google.android.apps.magazines:id/open_search_view_scrim",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        231
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 6,
    "resource_id": "com.google.android.apps.magazines:id/appbar",
    "scrollable": false,
    "selected": false,
    "size": "1080*231",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        84
      ],
      [
        1038,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      11,
      12
    ],
    "class": "android.widget.EditText",
    "clickable": true,
    "content_description": null,
    "editable": true,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 9,
    "resource_id": "com.google.android.apps.magazines:id/search_bar",
    "scrollable": false,
    "selected": false,
    "size": "996*126",
    "temp_id": 10,
    "text": "sustainable living",
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        84
      ],
      [
        179,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageButton",
    "clickable": true,
    "content_description": "Navigate up",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 10,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        179,
        116
      ],
      [
        889,
        178
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 10,
    "resource_id": "com.google.android.apps.magazines:id/open_search_bar_text_view",
    "scrollable": false,
    "selected": false,
    "size": "710*62",
    "temp_id": 12,
    "text": "sustainable living",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        231
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 8,
    "children": [
      14,
      23,
      24,
      36,
      37,
      53,
      68,
      84
    ],
    "class": "android.widget.ListView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 6,
    "resource_id": "com.google.android.apps.magazines:id/search_results_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*2169",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        231
      ],
      [
        1080,
        453
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      15,
      19,
      22
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*222",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        263
      ],
      [
        211,
        421
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      16
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 14,
    "resource_id": "com.google.android.apps.magazines:id/icon_frame",
    "scrollable": false,
    "selected": false,
    "size": "158*158",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        61,
        271
      ],
      [
        203,
        413
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      17
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 15,
    "resource_id": "com.google.android.apps.magazines:id/edition_icon_fixed_width",
    "scrollable": false,
    "selected": false,
    "size": "142*142",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        61,
        271
      ],
      [
        203,
        413
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 16,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "142*142",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        61,
        271
      ],
      [
        203,
        413
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 17,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "142*142",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        258,
        274
      ],
      [
        911,
        409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      20,
      21
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "653*135",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        258,
        274
      ],
      [
        911,
        353
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "653*79",
    "temp_id": 20,
    "text": "Sustainable Living News",
    "visible": true
  },
  {
    "bounds": [
      [
        258,
        353
      ],
      [
        911,
        409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "653*56",
    "temp_id": 21,
    "text": "Source",
    "visible": true
  },
  {
    "bounds": [
      [
        943,
        300
      ],
      [
        1027,
        384
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Follow",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 14,
    "resource_id": "com.google.android.apps.magazines:id/follow_button",
    "scrollable": false,
    "selected": false,
    "size": "84*84",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        453
      ],
      [
        1080,
        479
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*26",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        479
      ],
      [
        1080,
        1093
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      25,
      28
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*614",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        479
      ],
      [
        1080,
        655
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": "Sources",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 24,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*176",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        532
      ],
      [
        1080,
        602
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      27
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1027*70",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        532
      ],
      [
        1048,
        602
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 26,
    "resource_id": "com.google.android.apps.magazines:id/shelf_header_title",
    "scrollable": false,
    "selected": false,
    "size": "995*70",
    "temp_id": 27,
    "text": "Sources",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        655
      ],
      [
        1080,
        1040
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 24,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*385",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        655
      ],
      [
        1080,
        1040
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 28,
    "resource_id": "com.google.android.apps.magazines:id/carousel",
    "scrollable": false,
    "selected": false,
    "size": "1080*385",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        48,
        655
      ],
      [
        330,
        1040
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      31,
      35
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": "Sustainable Living News",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 29,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "282*385",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        48,
        655
      ],
      [
        330,
        937
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "282*282",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        56,
        663
      ],
      [
        322,
        929
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      33
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 31,
    "resource_id": "com.google.android.apps.magazines:id/edition_icon",
    "scrollable": false,
    "selected": false,
    "size": "266*266",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        56,
        663
      ],
      [
        322,
        929
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      34
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "266*266",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        56,
        663
      ],
      [
        322,
        929
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 33,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "266*266",
    "temp_id": 34,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        48,
        937
      ],
      [
        330,
        1040
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 30,
    "resource_id": "com.google.android.apps.magazines:id/source_name",
    "scrollable": false,
    "selected": false,
    "size": "282*103",
    "temp_id": 35,
    "text": "Sustainable Living News",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1093
      ],
      [
        1080,
        1119
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*26",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1151
      ],
      [
        1080,
        1556
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      38
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": "com.google.android.apps.magazines:id/card",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1151
      ],
      [
        1080,
        1556
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      39,
      50
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 37,
    "resource_id": "com.google.android.apps.magazines:id/card_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1198
      ],
      [
        1027,
        1429
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      40,
      47
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "974*231",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1198
      ],
      [
        796,
        1423
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      41,
      46
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "743*225",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1198
      ],
      [
        764,
        1238
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      45
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "711*40",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1199
      ],
      [
        90,
        1236
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 41,
    "resource_id": "com.google.android.apps.magazines:id/source_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1199
      ],
      [
        90,
        1236
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 42,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1199
      ],
      [
        90,
        1236
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 43,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        111,
        1198
      ],
      [
        764,
        1238
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "653*40",
    "temp_id": 45,
    "text": "WABE 90.1 FM",
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1254
      ],
      [
        764,
        1423
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 40,
    "resource_id": "com.google.android.apps.magazines:id/title",
    "scrollable": false,
    "selected": false,
    "size": "711*169",
    "temp_id": 46,
    "text": "MicroLife Institute promotes sustainable living through latest development \u2013 WABE",
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1198
      ],
      [
        1027,
        1429
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      48
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 47,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1198
      ],
      [
        1027,
        1429
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      49
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 47,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1198
      ],
      [
        1027,
        1429
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 48,
    "resource_id": "com.google.android.apps.magazines:id/image",
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 49,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1429
      ],
      [
        1080,
        1556
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      51,
      52
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1027*127",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1445
      ],
      [
        987,
        1540
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "6 hours ago",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 50,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "934*95",
    "temp_id": 51,
    "text": "6 hours ago",
    "visible": true
  },
  {
    "bounds": [
      [
        987,
        1445
      ],
      [
        1080,
        1540
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "More options",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 50,
    "resource_id": "com.google.android.apps.magazines:id/more_button",
    "scrollable": false,
    "selected": false,
    "size": "93*95",
    "temp_id": 52,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1556
      ],
      [
        1080,
        1961
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      54
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": "com.google.android.apps.magazines:id/card",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 53,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1556
      ],
      [
        1080,
        1961
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      55,
      65
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 53,
    "resource_id": "com.google.android.apps.magazines:id/card_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1603
      ],
      [
        1027,
        1834
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      56,
      62
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "974*231",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1603
      ],
      [
        796,
        1828
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      57,
      61
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "743*225",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1603
      ],
      [
        764,
        1643
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      58
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 56,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "711*40",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1604
      ],
      [
        127,
        1641
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      59
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": "TriplePundit",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 57,
    "resource_id": "com.google.android.apps.magazines:id/source_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "74*37",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1604
      ],
      [
        127,
        1641
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      60
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "74*37",
    "temp_id": 59,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1604
      ],
      [
        127,
        1641
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 59,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "74*37",
    "temp_id": 60,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1659
      ],
      [
        764,
        1828
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 56,
    "resource_id": "com.google.android.apps.magazines:id/title",
    "scrollable": false,
    "selected": false,
    "size": "711*169",
    "temp_id": 61,
    "text": "2024 Sustainable Living Challenge: Join Us in Making a Difference This Year",
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1603
      ],
      [
        1027,
        1834
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      63
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1603
      ],
      [
        1027,
        1834
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      64
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 62,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 63,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        1603
      ],
      [
        1027,
        1834
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 63,
    "resource_id": "com.google.android.apps.magazines:id/image",
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1834
      ],
      [
        1080,
        1961
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      66,
      67
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1027*127",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        1850
      ],
      [
        987,
        1945
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "6 days ago",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "934*95",
    "temp_id": 66,
    "text": "6 days ago",
    "visible": true
  },
  {
    "bounds": [
      [
        987,
        1850
      ],
      [
        1080,
        1945
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "More options",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 65,
    "resource_id": "com.google.android.apps.magazines:id/more_button",
    "scrollable": false,
    "selected": false,
    "size": "93*95",
    "temp_id": 67,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1961
      ],
      [
        1080,
        2366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      69
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": "com.google.android.apps.magazines:id/card",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 68,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1961
      ],
      [
        1080,
        2366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      70,
      81
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 68,
    "resource_id": "com.google.android.apps.magazines:id/card_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*405",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2008
      ],
      [
        1027,
        2239
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      71,
      78
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "974*231",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2008
      ],
      [
        796,
        2180
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      72,
      77
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 70,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "743*172",
    "temp_id": 71,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2008
      ],
      [
        764,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      73,
      76
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 71,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "711*40",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2009
      ],
      [
        90,
        2046
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      74
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 72,
    "resource_id": "com.google.android.apps.magazines:id/source_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 73,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2009
      ],
      [
        90,
        2046
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      75
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 73,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 74,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2009
      ],
      [
        90,
        2046
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 74,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 75,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        111,
        2008
      ],
      [
        764,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 72,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "653*40",
    "temp_id": 76,
    "text": "Blue & Green Tomorrow",
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2064
      ],
      [
        764,
        2180
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 71,
    "resource_id": "com.google.android.apps.magazines:id/title",
    "scrollable": false,
    "selected": false,
    "size": "711*116",
    "temp_id": 77,
    "text": "5 Tips for Creating a Sustainable Living Space",
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        2008
      ],
      [
        1027,
        2239
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      79
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 70,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 78,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        2008
      ],
      [
        1027,
        2239
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      80
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 78,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 79,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        796,
        2008
      ],
      [
        1027,
        2239
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 79,
    "resource_id": "com.google.android.apps.magazines:id/image",
    "scrollable": false,
    "selected": false,
    "size": "231*231",
    "temp_id": 80,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2239
      ],
      [
        1080,
        2366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      82,
      83
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1027*127",
    "temp_id": 81,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        53,
        2255
      ],
      [
        987,
        2350
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "6 days ago",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 81,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "934*95",
    "temp_id": 82,
    "text": "6 days ago",
    "visible": true
  },
  {
    "bounds": [
      [
        987,
        2255
      ],
      [
        1080,
        2350
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "More options",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 81,
    "resource_id": "com.google.android.apps.magazines:id/more_button",
    "scrollable": false,
    "selected": false,
    "size": "93*95",
    "temp_id": 83,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2366
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      85
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 13,
    "resource_id": "com.google.android.apps.magazines:id/card",
    "scrollable": false,
    "selected": false,
    "size": "1080*34",
    "temp_id": 84,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2366
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      86,
      96
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 84,
    "resource_id": "com.google.android.apps.magazines:id/card_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*34",
    "temp_id": 85,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2413
      ],
      [
        1027,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      87,
      93
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 85,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "974*-13",
    "temp_id": 86,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2413
      ],
      [
        796,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      88,
      92
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 86,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "743*-13",
    "temp_id": 87,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2413
      ],
      [
        764,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      89
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 87,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "711*-13",
    "temp_id": 88,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2414
      ],
      [
        316,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      90
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": "Yahoo Finance",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 88,
    "resource_id": "com.google.android.apps.magazines:id/source_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "263*-14",
    "temp_id": 89,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2414
      ],
      [
        316,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      91
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 89,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "263*-14",
    "temp_id": 90,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2414
      ],
      [
        316,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 90,
    "resource_id": "com.google.android.apps.magazines:id/rect_icon",
    "scrollable": false,
    "selected": false,
    "size": "263*-14",
    "temp_id": 91,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2469
      ],
      [
        764,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 87,
    "resource_id": "com.google.android.apps.magazines:id/title",
    "scrollable": false,
    "selected": false,
    "size": "711*-69",
    "temp_id": 92,
    "text": "Hydrofarm Showcases Sustainable Indoor Gardening Solutions on 'The Balancing Act'",
    "visible": false
  },
  {
    "bounds": [
      [
        796,
        2413
      ],
      [
        1027,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      94
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 86,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*-13",
    "temp_id": 93,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        796,
        2413
      ],
      [
        1027,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      95
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 93,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*-13",
    "temp_id": 94,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        796,
        2413
      ],
      [
        1027,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 94,
    "resource_id": "com.google.android.apps.magazines:id/image",
    "scrollable": false,
    "selected": false,
    "size": "231*-13",
    "temp_id": 95,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2644
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      97,
      98
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 85,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1027*-244",
    "temp_id": 96,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        53,
        2660
      ],
      [
        987,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "5 days ago",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 96,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "934*-260",
    "temp_id": 97,
    "text": "5 days ago",
    "visible": false
  },
  {
    "bounds": [
      [
        987,
        2660
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "More options",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 96,
    "resource_id": "com.google.android.apps.magazines:id/more_button",
    "scrollable": false,
    "selected": false,
    "size": "93*-260",
    "temp_id": 98,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2274
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.magazines",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 99,
    "text": null,
    "visible": false
  }
]
