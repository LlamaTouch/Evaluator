[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      74
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      73
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 9,
    "children": [
      7,
      8,
      9,
      10,
      11,
      12,
      13,
      69,
      72
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 10,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": "com.google.android.apps.maps:id/fullscreen_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      16
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      17,
      27
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar",
    "scrollable": false,
    "selected": false,
    "size": "1080*211",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*148",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      20,
      21,
      24
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/toolbar",
    "scrollable": false,
    "selected": false,
    "size": "1080*148",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1059,
        63
      ],
      [
        1059,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/end_section",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 20,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        21,
        63
      ],
      [
        168,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/start_section",
    "scrollable": false,
    "selected": false,
    "size": "147*148",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        74
      ],
      [
        147,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      23
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Navigate up",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/nav_button",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        74
      ],
      [
        147,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar_button_icon",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        168,
        63
      ],
      [
        912,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      25
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/title_frame",
    "scrollable": false,
    "selected": false,
    "size": "744*148",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        364,
        74
      ],
      [
        716,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 24,
    "resource_id": "com.google.android.apps.maps:id/title_section",
    "scrollable": false,
    "selected": false,
    "size": "352*126",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        364,
        103
      ],
      [
        716,
        171
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 25,
    "resource_id": "com.google.android.apps.maps:id/title",
    "scrollable": false,
    "selected": false,
    "size": "352*68",
    "temp_id": 26,
    "text": "Personal content",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      28
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar_fullscreen_content_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 27,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 29,
    "resource_id": "android:id/list_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 9,
    "children": [
      32,
      35,
      41,
      47,
      50,
      54,
      57,
      61,
      65
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        223
      ],
      [
        1080,
        316
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      33
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        223
      ],
      [
        1038,
        316
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      34
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        244
      ],
      [
        1038,
        295
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 34,
    "text": "Your Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        316
      ],
      [
        1080,
        508
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      36,
      39
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*192",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        316
      ],
      [
        874,
        508
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      37,
      38
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*192",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        358
      ],
      [
        335,
        415
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "293*57",
    "temp_id": 37,
    "text": "Timeline emails",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        415
      ],
      [
        759,
        466
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "717*51",
    "temp_id": 38,
    "text": "Get highlights of your Timeline in your inbox",
    "visible": true
  },
  {
    "bounds": [
      [
        874,
        316
      ],
      [
        1038,
        508
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      40
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": "android:id/widget_frame",
    "scrollable": false,
    "selected": false,
    "size": "164*192",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        916,
        376
      ],
      [
        1038,
        447
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Switch",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 39,
    "resource_id": "com.google.android.apps.maps:id/switchWidget",
    "scrollable": false,
    "selected": false,
    "size": "122*71",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        508
      ],
      [
        1080,
        700
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      45
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*192",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        508
      ],
      [
        874,
        700
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      43,
      44
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*192",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        550
      ],
      [
        319,
        607
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "277*57",
    "temp_id": 43,
    "text": "Google Photos",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        607
      ],
      [
        653,
        658
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "611*51",
    "temp_id": 44,
    "text": "Show your Google Photos in Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        874,
        508
      ],
      [
        1038,
        700
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      46
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": "android:id/widget_frame",
    "scrollable": false,
    "selected": false,
    "size": "164*192",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        916,
        568
      ],
      [
        1038,
        639
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Switch",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 45,
    "resource_id": "com.google.android.apps.maps:id/switchWidget",
    "scrollable": false,
    "selected": false,
    "size": "122*71",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        745
      ],
      [
        1080,
        838
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      48
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 47,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        745
      ],
      [
        1038,
        838
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      49
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 47,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        766
      ],
      [
        1038,
        817
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 48,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 49,
    "text": "App history",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        838
      ],
      [
        1080,
        1073
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      51
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        838
      ],
      [
        1038,
        1073
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      52,
      53
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 50,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        880
      ],
      [
        507,
        937
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "465*57",
    "temp_id": 52,
    "text": "Web & App Activity is off\u00a0",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        937
      ],
      [
        1038,
        1031
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 53,
    "text": "Allow features to work properly like Timeline and search suggestions",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1115
      ],
      [
        1080,
        1208
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      55
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1115
      ],
      [
        1038,
        1208
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1136
      ],
      [
        1038,
        1187
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 56,
    "text": "Location settings",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1208
      ],
      [
        1080,
        1443
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      58
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1208
      ],
      [
        1038,
        1443
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      59,
      60
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 57,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1250
      ],
      [
        304,
        1307
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "262*57",
    "temp_id": 59,
    "text": "Location is on",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1307
      ],
      [
        1038,
        1401
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 60,
    "text": "Let this app know your location for things like directions, navigation and search",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1443
      ],
      [
        1080,
        1678
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      62
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 61,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1443
      ],
      [
        1038,
        1678
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      63,
      64
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1485
      ],
      [
        300,
        1542
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "258*57",
    "temp_id": 63,
    "text": "Timeline is on",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1542
      ],
      [
        1038,
        1636
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 64,
    "text": "Rediscover the places you've been and the routes you've traveled",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1678
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      66
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*114",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1678
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      67,
      68
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*114",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1720
      ],
      [
        476,
        1777
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 66,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "434*57",
    "temp_id": 67,
    "text": "Delete all Timeline data",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1777
      ],
      [
        911,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 66,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "869*15",
    "temp_id": 68,
    "text": "Permanently delete visits and routes from this device",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      70
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      71
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 71,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 73,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 74,
    "text": null,
    "visible": false
  }
]
