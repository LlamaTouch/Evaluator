[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      1,
      52,
      53
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 2,
    "resource_id": "com.google.android.apps.photos:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      7
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 4,
    "resource_id": "com.google.android.apps.photos:id/touch_capture_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 5,
    "resource_id": "com.google.android.apps.photos:id/photo_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "androidx.drawerlayout.widget.DrawerLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 5,
    "resource_id": "com.google.android.apps.photos:id/drawer_layout",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      9
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 7,
    "resource_id": "com.google.android.apps.photos:id/main_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      10,
      25,
      42
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 8,
    "resource_id": "com.google.android.apps.photos:id/toolbar_parent",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 9,
    "resource_id": "com.google.android.apps.photos:id/touch_capture_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      12,
      20,
      24
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 10,
    "resource_id": "com.google.android.apps.photos:id/all_photos_coordinator",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      13
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 11,
    "resource_id": "com.google.android.apps.photos:id/fragment_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      14,
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 12,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 13,
    "resource_id": "com.google.android.apps.photos:id/fragment_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      16
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 14,
    "resource_id": "com.google.android.apps.photos:id/fragment_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      17
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 15,
    "resource_id": "com.google.android.apps.photos:id/photos_photogrid_date_scrubber_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 16,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1645
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 17,
    "resource_id": "com.google.android.apps.photos:id/recycler_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1645",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 13,
    "resource_id": "com.google.android.apps.photos:id/empty_view_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      21,
      22,
      23
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 11,
    "resource_id": "com.google.android.apps.photos:id/all_photos_empty_state_layout",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        251,
        638
      ],
      [
        829,
        843
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": "No photos",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "578*205",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        943
      ],
      [
        907,
        1075
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*132",
    "temp_id": 22,
    "text": "No photos",
    "visible": true
  },
  {
    "bounds": [
      [
        172,
        1075
      ],
      [
        907,
        1237
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "735*162",
    "temp_id": 23,
    "text": "Take a picture. Photos & videos appear here.",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1876
      ],
      [
        1038,
        1876
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 11,
    "resource_id": "com.google.android.apps.photos:id/hats_container",
    "scrollable": false,
    "selected": false,
    "size": "996*0",
    "temp_id": 24,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 9,
    "resource_id": "com.google.android.apps.photos:id/scrolling_toolbar_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*210",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      27,
      28
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 25,
    "resource_id": "com.google.android.apps.photos:id/toolbar_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*210",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 26,
    "resource_id": "com.google.android.apps.photos:id/notification_bar_spacer",
    "scrollable": false,
    "selected": false,
    "size": "1080*63",
    "temp_id": 27,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      29,
      30,
      35
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 26,
    "resource_id": "com.google.android.apps.photos:id/toolbar",
    "scrollable": false,
    "selected": false,
    "size": "1080*147",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        147,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageButton",
    "clickable": true,
    "content_description": "Printing",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "147*147",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        368,
        63
      ],
      [
        712,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      31,
      34
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "344*147",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        368,
        104
      ],
      [
        712,
        169
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      32,
      33
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": "Google Photos",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 30,
    "resource_id": "com.google.android.apps.photos:id/product_lockup_view",
    "scrollable": false,
    "selected": false,
    "size": "344*65",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        368,
        111
      ],
      [
        546,
        169
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 31,
    "resource_id": "com.google.android.apps.photos:id/logo",
    "scrollable": false,
    "selected": false,
    "size": "178*58",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        556,
        104
      ],
      [
        712,
        167
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 31,
    "resource_id": "com.google.android.apps.photos:id/product_name",
    "scrollable": false,
    "selected": false,
    "size": "156*63",
    "temp_id": 33,
    "text": "Photos",
    "visible": true
  },
  {
    "bounds": [
      [
        540,
        143
      ],
      [
        540,
        186
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 30,
    "resource_id": "com.google.android.apps.photos:id/message_text_view",
    "scrollable": false,
    "selected": false,
    "size": "0*43",
    "temp_id": 34,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        933,
        63
      ],
      [
        1080,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      36
    ],
    "class": "android.support.v7.widget.LinearLayoutCompat",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "147*147",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        933,
        73
      ],
      [
        1080,
        199
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      37
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Signed in as Ian agentian03@gmail.com\nBackup is off.\nAccount and settings.",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 35,
    "resource_id": "com.google.android.apps.photos:id/selected_account_disc",
    "scrollable": false,
    "selected": false,
    "size": "147*126",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        933,
        73
      ],
      [
        1059,
        199
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      38,
      39,
      40
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 36,
    "resource_id": "com.google.android.apps.photos:id/og_selected_account_disc_apd",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        938,
        78
      ],
      [
        1054,
        194
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 37,
    "resource_id": "com.google.android.apps.photos:id/og_apd_internal_image_view",
    "scrollable": false,
    "selected": false,
    "size": "116*116",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        938,
        78
      ],
      [
        1054,
        194
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 37,
    "resource_id": "com.google.android.apps.photos:id/og_apd_ring_view",
    "scrollable": false,
    "selected": false,
    "size": "116*116",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1004,
        144
      ],
      [
        1051,
        191
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      41
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 37,
    "resource_id": "com.google.android.apps.photos:id/badge_wrapper",
    "scrollable": false,
    "selected": false,
    "size": "47*47",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1009,
        149
      ],
      [
        1046,
        186
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 40,
    "resource_id": "com.google.android.apps.photos:id/og_apd_drawable_badge",
    "scrollable": false,
    "selected": false,
    "size": "37*37",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1632
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 9,
    "resource_id": "com.google.android.apps.photos:id/tab_bar",
    "scrollable": false,
    "selected": false,
    "size": "1080*286",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1632
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 42,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*286",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1632
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      45,
      46,
      51
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 43,
    "resource_id": "com.google.android.apps.photos:id/tab_layout",
    "scrollable": false,
    "selected": false,
    "size": "1080*286",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1632
      ],
      [
        1080,
        1645
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 44,
    "resource_id": "com.google.android.apps.photos:id/tab_bar_top_shadow",
    "scrollable": false,
    "selected": false,
    "size": "1080*13",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1645
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      47,
      48,
      49,
      50
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*147",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1645
      ],
      [
        270,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 46,
    "resource_id": "com.google.android.apps.photos:id/tab_photos",
    "scrollable": false,
    "selected": true,
    "size": "270*147",
    "temp_id": 47,
    "text": "Photos",
    "visible": true
  },
  {
    "bounds": [
      [
        270,
        1645
      ],
      [
        540,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.photos",
    "parent": 46,
    "resource_id": "com.google.android.apps.photos:id/search_destination",
    "scrollable": false,
    "selected": false,
    "size": "270*147",
    "temp_id": 48,
    "text": "Search",
    "visible": true
  },
  {
    "bounds": [
      [
        540,
        1645
      ],
      [
        810,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 46,
    "resource_id": "com.google.android.apps.photos:id/tab_sharing",
    "scrollable": false,
    "selected": false,
    "size": "270*147",
    "temp_id": 49,
    "text": "Sharing",
    "visible": true
  },
  {
    "bounds": [
      [
        810,
        1645
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 46,
    "resource_id": "com.google.android.apps.photos:id/tab_library",
    "scrollable": false,
    "selected": false,
    "size": "270*147",
    "temp_id": 50,
    "text": "Library",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 44,
    "resource_id": "com.google.android.apps.photos:id/fill_under_navigation_bar",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 51,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 0,
    "resource_id": "android:id/statusBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*63",
    "temp_id": 52,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.photos",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 53,
    "text": null,
    "visible": false
  }
]
