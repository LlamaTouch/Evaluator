[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      71
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      70
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 10,
    "children": [
      7,
      8,
      9,
      10,
      13,
      14,
      16,
      17,
      18,
      69
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        661
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1071*126",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        661
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      12
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 10,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1071*126",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        535
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 11,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1071*0",
    "temp_id": 12,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 13,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/map_frame",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      20
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/fullscreen_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      21
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      23
    ],
    "class": "android.webkit.WebView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      24
    ],
    "class": "android.webkit.WebView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": true,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 23,
    "text": "Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      25
    ],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 23,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 24,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 24,
    "resource_id": "yDmH0d",
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 25,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      27
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 26,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      28
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 27,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 28,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 29,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      31,
      61,
      64
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 29,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 30,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*336",
    "temp_id": 31,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      33,
      53,
      60
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*273",
    "temp_id": 32,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1084,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      34,
      36,
      37,
      39
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*147",
    "temp_id": 33,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        196
      ],
      [
        1084,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      35
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*14",
    "temp_id": 34,
    "text": "Back",
    "visible": false
  },
  {
    "bounds": [
      [
        7,
        70
      ],
      [
        139,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 34,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 35,
    "text": "Back",
    "visible": false
  },
  {
    "bounds": [
      [
        126,
        105
      ],
      [
        958,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*63",
    "temp_id": 36,
    "text": "Timeline",
    "visible": false
  },
  {
    "bounds": [
      [
        805,
        70
      ],
      [
        937,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      38
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 37,
    "text": "Backup disabled.",
    "visible": false
  },
  {
    "bounds": [
      [
        805,
        70
      ],
      [
        937,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 38,
    "text": "Backup disabled.",
    "visible": false
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      40
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 39,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      41,
      43
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 40,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      42
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 41,
    "text": "More options",
    "visible": false
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 42,
    "text": "More options",
    "visible": false
  },
  {
    "bounds": [
      [
        498,
        196
      ],
      [
        1071,
        1170
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*974",
    "temp_id": 43,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        196
      ],
      [
        1071,
        1170
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 8,
    "children": [
      45,
      46,
      47,
      48,
      49,
      50,
      51,
      52
    ],
    "class": "android.widget.ListView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 43,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*974",
    "temp_id": 44,
    "text": "Options list",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        217
      ],
      [
        1071,
        349
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*132",
    "temp_id": 45,
    "text": "About Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        343
      ],
      [
        1071,
        475
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*132",
    "temp_id": 46,
    "text": "Settings and privacy",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        469
      ],
      [
        1071,
        601
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*132",
    "temp_id": 47,
    "text": "Help",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        595
      ],
      [
        1071,
        727
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*132",
    "temp_id": 48,
    "text": "Send feedback",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        742
      ],
      [
        1071,
        750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*8",
    "temp_id": 49,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        766
      ],
      [
        1071,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*131",
    "temp_id": 50,
    "text": "Refresh",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        892
      ],
      [
        1071,
        1023
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*131",
    "temp_id": 51,
    "text": "Delete day",
    "visible": true
  },
  {
    "bounds": [
      [
        498,
        1018
      ],
      [
        1071,
        1149
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.MenuItem",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "573*131",
    "temp_id": 52,
    "text": "Add to Home screen",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 6,
    "children": [
      54,
      55,
      56,
      57,
      58,
      59
    ],
    "class": "android.widget.TabWidget",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*126",
    "temp_id": 53,
    "text": "",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        154,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab1",
    "scrollable": false,
    "selected": true,
    "size": "154*126",
    "temp_id": 54,
    "text": "Day",
    "visible": false
  },
  {
    "bounds": [
      [
        149,
        210
      ],
      [
        325,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab5",
    "scrollable": false,
    "selected": false,
    "size": "176*126",
    "temp_id": 55,
    "text": "Trips",
    "visible": false
  },
  {
    "bounds": [
      [
        320,
        210
      ],
      [
        546,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab6",
    "scrollable": false,
    "selected": false,
    "size": "226*126",
    "temp_id": 56,
    "text": "Insights",
    "visible": false
  },
  {
    "bounds": [
      [
        543,
        210
      ],
      [
        745,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab2",
    "scrollable": false,
    "selected": false,
    "size": "202*126",
    "temp_id": 57,
    "text": "Places",
    "visible": false
  },
  {
    "bounds": [
      [
        742,
        210
      ],
      [
        931,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab3",
    "scrollable": false,
    "selected": false,
    "size": "189*126",
    "temp_id": 58,
    "text": "Cities",
    "visible": false
  },
  {
    "bounds": [
      [
        926,
        210
      ],
      [
        1120,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": "tab4",
    "scrollable": false,
    "selected": false,
    "size": "194*126",
    "temp_id": 59,
    "text": "World",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        336
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*0",
    "temp_id": 60,
    "text": "",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        336
      ],
      [
        1084,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      62,
      63
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*561",
    "temp_id": 61,
    "text": "Timeline is on Past visits layer is off",
    "visible": false
  },
  {
    "bounds": [
      [
        910,
        364
      ],
      [
        1042,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 62,
    "text": "Timeline is on",
    "visible": false
  },
  {
    "bounds": [
      [
        910,
        748
      ],
      [
        1042,
        876
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*128",
    "temp_id": 63,
    "text": "Past visits layer is off",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        895
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      65,
      66,
      67,
      68
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*898",
    "temp_id": 64,
    "text": "Previous day Today No visits for this day Edit",
    "visible": false
  },
  {
    "bounds": [
      [
        -1063,
        947
      ],
      [
        -931,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*129",
    "temp_id": 65,
    "text": "Previous day",
    "visible": false
  },
  {
    "bounds": [
      [
        -149,
        947
      ],
      [
        -21,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "128*129",
    "temp_id": 66,
    "text": "Next day",
    "visible": false
  },
  {
    "bounds": [
      [
        18,
        947
      ],
      [
        147,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "129*129",
    "temp_id": 67,
    "text": "Previous day",
    "visible": false
  },
  {
    "bounds": [
      [
        897,
        1609
      ],
      [
        1050,
        1761
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "153*152",
    "temp_id": 68,
    "text": "Edit",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 70,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 71,
    "text": null,
    "visible": false
  }
]
