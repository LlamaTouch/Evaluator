[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      149
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      148
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 15,
    "children": [
      7,
      8,
      9,
      11,
      12,
      13,
      35,
      80,
      88,
      100,
      101,
      135,
      136,
      137,
      140
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/map_frame",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 9,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        226
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        226
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      15,
      16
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        226
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        226
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      17
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        15,
        60
      ],
      [
        1065,
        226
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1050*166",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      20
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      21
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      22,
      25,
      29,
      34
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": "com.google.android.apps.maps:id/mod_search_omnibox_layout",
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        789,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      23,
      24
    ],
    "class": "android.widget.EditText",
    "clickable": true,
    "content_description": "Search here",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_text_box",
    "scrollable": false,
    "selected": false,
    "size": "758*126",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        62,
        110
      ],
      [
        136,
        184
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "74*74",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        162,
        84
      ],
      [
        789,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "627*126",
    "temp_id": 24,
    "text": "Search here",
    "visible": true
  },
  {
    "bounds": [
      [
        789,
        84
      ],
      [
        915,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        789,
        84
      ],
      [
        915,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      27
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        789,
        84
      ],
      [
        915,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      28
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 27,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        789,
        84
      ],
      [
        915,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        915,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_one_google_account_disc",
    "scrollable": false,
    "selected": false,
    "size": "134*126",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        915,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Signed in as Ian agentian03@gmail.com\nAccount and settings.",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 29,
    "resource_id": "com.google.android.apps.maps:id/selected_account_disc",
    "scrollable": false,
    "selected": false,
    "size": "134*126",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        915,
        84
      ],
      [
        1041,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      32,
      33
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": "com.google.android.apps.maps:id/og_selected_account_disc_apd",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        923,
        92
      ],
      [
        923,
        92
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": "com.google.android.apps.maps:id/ring_wrapper",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 32,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        923,
        92
      ],
      [
        1033,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": "com.google.android.apps.maps:id/og_apd_internal_image_view",
    "scrollable": false,
    "selected": false,
    "size": "110*110",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        915,
        147
      ],
      [
        915,
        147
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_live_view_entry_layout",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 34,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        226
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      36
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1566",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        226
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      37
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": "com.google.android.apps.maps:id/explore_tab_home_bottom_sheet",
    "scrollable": true,
    "selected": false,
    "size": "1080*1566",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1219
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      38,
      77
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*573",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1219
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      39,
      49
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": "Explore this area",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": "com.google.android.apps.maps:id/scrollable_card_stream_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*573",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1219
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      40
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*147",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1240
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      41
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1240
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      42
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1240
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1240
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "com.google.android.apps.maps:id/explore_tab_home_title_card",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1240
      ],
      [
        1080,
        1366
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      45,
      48
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 43,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1276
      ],
      [
        1080,
        1361
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      46
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*85",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1276
      ],
      [
        1028,
        1361
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      47
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 45,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*85",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1276
      ],
      [
        1028,
        1361
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*85",
    "temp_id": 47,
    "text": "Latest in the area",
    "visible": true
  },
  {
    "bounds": [
      [
        1080,
        1318
      ],
      [
        1080,
        1318
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 48,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1366
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      50
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*426",
    "temp_id": 49,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1366
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      51
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 49,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*426",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1366
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      52
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 50,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*426",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1366
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      53,
      64,
      67,
      73
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": "Post number 1, Posted a week ago",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*426",
    "temp_id": 52,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1387
      ],
      [
        1080,
        1528
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      54,
      62
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 52,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*141",
    "temp_id": 53,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1387
      ],
      [
        860,
        1528
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      55,
      58
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "860*141",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1415
      ],
      [
        157,
        1499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "105*84",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1415
      ],
      [
        136,
        1499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      57
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "84*84",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1415
      ],
      [
        136,
        1499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 56,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "84*84",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        1408
      ],
      [
        829,
        1507
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      59,
      60
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "672*99",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        1408
      ],
      [
        457,
        1464
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "com.google.android.apps.maps:id/textbox",
    "scrollable": false,
    "selected": false,
    "size": "300*56",
    "temp_id": 59,
    "text": "Ricardo Castelan",
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        1464
      ],
      [
        829,
        1507
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      61
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "672*43",
    "temp_id": 60,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        1464
      ],
      [
        829,
        1507
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 60,
    "resource_id": "com.google.android.apps.maps:id/textbox",
    "scrollable": false,
    "selected": false,
    "size": "672*43",
    "temp_id": 61,
    "text": "Local Guide \u00b7 2 photos",
    "visible": true
  },
  {
    "bounds": [
      [
        860,
        1394
      ],
      [
        1080,
        1520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      63
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "220*126",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        860,
        1394
      ],
      [
        1080,
        1520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "220*126",
    "temp_id": 63,
    "text": "Follow",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1528
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      65
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 52,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*264",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1538
      ],
      [
        1028,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      66
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": "Photo of Balneario Las Lumbreras",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*254",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        52,
        1538
      ],
      [
        1028,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*254",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2326
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      68,
      69,
      72
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 52,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-534",
    "temp_id": 67,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        52,
        2327
      ],
      [
        795,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 67,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "743*-535",
    "temp_id": 68,
    "text": "a week ago",
    "visible": false
  },
  {
    "bounds": [
      [
        795,
        2326
      ],
      [
        933,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      70,
      71
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Photo of Balneario Las Lumbreras by Ricardo Castelan, 199 people have liked this photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 67,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "138*-534",
    "temp_id": 69,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        795,
        2362
      ],
      [
        858,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "63*-570",
    "temp_id": 70,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        858,
        2363
      ],
      [
        933,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "75*-571",
    "temp_id": 71,
    "text": "199",
    "visible": false
  },
  {
    "bounds": [
      [
        933,
        2326
      ],
      [
        1059,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageButton",
    "clickable": true,
    "content_description": "More options for post by Ricardo Castelan",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 67,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-534",
    "temp_id": 72,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        52,
        2452
      ],
      [
        1028,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      74
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 52,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*-660",
    "temp_id": 73,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        52,
        2452
      ],
      [
        1028,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      75,
      76
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 73,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "976*-660",
    "temp_id": 74,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        94,
        2483
      ],
      [
        986,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 74,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "892*-691",
    "temp_id": 75,
    "text": "Balneario Las Lumbreras",
    "visible": false
  },
  {
    "bounds": [
      [
        94,
        2539
      ],
      [
        986,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 74,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "892*-747",
    "temp_id": 76,
    "text": "4.1 stars  \u2022  Water park  \u2022  Ajacuba",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1219
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      78
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*573",
    "temp_id": 77,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        613,
        2394
      ],
      [
        1067,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      79
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "454*-602",
    "temp_id": 78,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        645,
        2426
      ],
      [
        1036,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Add a post",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 78,
    "resource_id": "com.google.android.apps.maps:id/terra_floating_action_button_view_model_impl",
    "scrollable": false,
    "selected": false,
    "size": "391*-634",
    "temp_id": 79,
    "text": "Add a post",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        226
      ],
      [
        1080,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      81
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 80,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        226
      ],
      [
        1080,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      82
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 81,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        226
      ],
      [
        1080,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      83
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 81,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1049*126",
    "temp_id": 82,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        226
      ],
      [
        1080,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      84,
      85,
      86,
      87
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 82,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1049*126",
    "temp_id": 83,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        226
      ],
      [
        371,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Search for Restaurants",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 83,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "340*126",
    "temp_id": 84,
    "text": "Restaurants",
    "visible": true
  },
  {
    "bounds": [
      [
        386,
        226
      ],
      [
        586,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Search for Gas",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 83,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "200*126",
    "temp_id": 85,
    "text": "Gas",
    "visible": true
  },
  {
    "bounds": [
      [
        601,
        226
      ],
      [
        904,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Search for Groceries",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 83,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "303*126",
    "temp_id": 86,
    "text": "Groceries",
    "visible": true
  },
  {
    "bounds": [
      [
        919,
        226
      ],
      [
        1080,
        352
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Search for Hotels",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 83,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "161*126",
    "temp_id": 87,
    "text": "Hotels",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        363
      ],
      [
        1080,
        651
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      89
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*288",
    "temp_id": 88,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        363
      ],
      [
        1080,
        651
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      90
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 88,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*288",
    "temp_id": 89,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        363
      ],
      [
        1080,
        520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      91
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 89,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 90,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        363
      ],
      [
        1080,
        520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      92
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 90,
    "resource_id": "com.google.android.apps.maps:id/layers_fab_button",
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 91,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1080,
        520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      93
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 91,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 92,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1080,
        520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      94
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 92,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 93,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1080,
        520
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      95
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Layers",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 93,
    "resource_id": "com.google.android.apps.maps:id/layers_fab",
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 94,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1049,
        499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      96,
      98
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 94,
    "resource_id": "com.google.android.apps.maps:id/fab_icon",
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 95,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1049,
        499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      97
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 96,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1049,
        499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 96,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 97,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1049,
        499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      99
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 98,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        378
      ],
      [
        1049,
        499
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 98,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 99,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 100,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1624
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      102
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/footer_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*168",
    "temp_id": 101,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1624
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      103
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 101,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*168",
    "temp_id": 102,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1624
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      104
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 102,
    "resource_id": "com.google.android.apps.maps:id/bottom_nav",
    "scrollable": false,
    "selected": false,
    "size": "1080*168",
    "temp_id": 103,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1624
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      105,
      111,
      117,
      123,
      129
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 103,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*168",
    "temp_id": 104,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1624
      ],
      [
        216,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      106,
      109
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": "Explore",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 104,
    "resource_id": "com.google.android.apps.maps:id/explore_tab_strip_button",
    "scrollable": false,
    "selected": true,
    "size": "216*168",
    "temp_id": 105,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        24,
        1635
      ],
      [
        192,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      107,
      108
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 105,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_container",
    "scrollable": false,
    "selected": true,
    "size": "168*84",
    "temp_id": 106,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        24,
        1635
      ],
      [
        192,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 106,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_active_indicator_view",
    "scrollable": false,
    "selected": true,
    "size": "168*84",
    "temp_id": 107,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        76,
        1645
      ],
      [
        139,
        1708
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 106,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_view",
    "scrollable": false,
    "selected": true,
    "size": "63*63",
    "temp_id": 108,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        1724
      ],
      [
        166,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      110
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 105,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_labels_group",
    "scrollable": false,
    "selected": true,
    "size": "116*68",
    "temp_id": 109,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        1724
      ],
      [
        166,
        1774
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 109,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_large_label_view",
    "scrollable": false,
    "selected": true,
    "size": "116*50",
    "temp_id": 110,
    "text": "Explore",
    "visible": true
  },
  {
    "bounds": [
      [
        216,
        1624
      ],
      [
        432,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      112,
      115
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Go",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 104,
    "resource_id": "com.google.android.apps.maps:id/transportation_tab_strip_button",
    "scrollable": false,
    "selected": false,
    "size": "216*168",
    "temp_id": 111,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        240,
        1635
      ],
      [
        408,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      113,
      114
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 111,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "168*84",
    "temp_id": 112,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        290,
        1635
      ],
      [
        358,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 112,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_active_indicator_view",
    "scrollable": false,
    "selected": false,
    "size": "68*84",
    "temp_id": 113,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        292,
        1645
      ],
      [
        355,
        1708
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 112,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_view",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 114,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        302,
        1724
      ],
      [
        346,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      116
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 111,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_labels_group",
    "scrollable": false,
    "selected": false,
    "size": "44*68",
    "temp_id": 115,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        302,
        1724
      ],
      [
        346,
        1774
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 115,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_small_label_view",
    "scrollable": false,
    "selected": false,
    "size": "44*50",
    "temp_id": 116,
    "text": "Go",
    "visible": true
  },
  {
    "bounds": [
      [
        432,
        1624
      ],
      [
        648,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      118,
      121
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Saved",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 104,
    "resource_id": "com.google.android.apps.maps:id/saved_tab_strip_button",
    "scrollable": false,
    "selected": false,
    "size": "216*168",
    "temp_id": 117,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        456,
        1635
      ],
      [
        624,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      119,
      120
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 117,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "168*84",
    "temp_id": 118,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        506,
        1635
      ],
      [
        574,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 118,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_active_indicator_view",
    "scrollable": false,
    "selected": false,
    "size": "68*84",
    "temp_id": 119,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        508,
        1645
      ],
      [
        571,
        1708
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 118,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_view",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 120,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        492,
        1724
      ],
      [
        588,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      122
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 117,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_labels_group",
    "scrollable": false,
    "selected": false,
    "size": "96*68",
    "temp_id": 121,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        492,
        1724
      ],
      [
        588,
        1774
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 121,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_small_label_view",
    "scrollable": false,
    "selected": false,
    "size": "96*50",
    "temp_id": 122,
    "text": "Saved",
    "visible": true
  },
  {
    "bounds": [
      [
        648,
        1624
      ],
      [
        864,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      124,
      127
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Contribute",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 104,
    "resource_id": "com.google.android.apps.maps:id/contribute_tab_strip_button",
    "scrollable": false,
    "selected": false,
    "size": "216*168",
    "temp_id": 123,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        672,
        1635
      ],
      [
        840,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      125,
      126
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 123,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "168*84",
    "temp_id": 124,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        722,
        1635
      ],
      [
        790,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 124,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_active_indicator_view",
    "scrollable": false,
    "selected": false,
    "size": "68*84",
    "temp_id": 125,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        724,
        1645
      ],
      [
        787,
        1708
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 124,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_view",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 126,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        673,
        1724
      ],
      [
        839,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      128
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 123,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_labels_group",
    "scrollable": false,
    "selected": false,
    "size": "166*68",
    "temp_id": 127,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        673,
        1724
      ],
      [
        839,
        1774
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 127,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_small_label_view",
    "scrollable": false,
    "selected": false,
    "size": "166*50",
    "temp_id": 128,
    "text": "Contribute",
    "visible": true
  },
  {
    "bounds": [
      [
        864,
        1624
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      130,
      133
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Updates",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 104,
    "resource_id": "com.google.android.apps.maps:id/updates_tab_strip_button",
    "scrollable": false,
    "selected": false,
    "size": "216*168",
    "temp_id": 129,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        888,
        1635
      ],
      [
        1056,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      131,
      132
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 129,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_container",
    "scrollable": false,
    "selected": false,
    "size": "168*84",
    "temp_id": 130,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        938,
        1635
      ],
      [
        1006,
        1719
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 130,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_active_indicator_view",
    "scrollable": false,
    "selected": false,
    "size": "68*84",
    "temp_id": 131,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        940,
        1645
      ],
      [
        1003,
        1708
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 130,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_icon_view",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 132,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        907,
        1724
      ],
      [
        1036,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      134
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 129,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_labels_group",
    "scrollable": false,
    "selected": false,
    "size": "129*68",
    "temp_id": 133,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        907,
        1724
      ],
      [
        1036,
        1774
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 133,
    "resource_id": "com.google.android.apps.maps:id/navigation_bar_item_small_label_view",
    "scrollable": false,
    "selected": false,
    "size": "129*50",
    "temp_id": 134,
    "text": "Updates",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1127
      ],
      [
        215,
        1193
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/watermark_image",
    "scrollable": false,
    "selected": false,
    "size": "173*66",
    "temp_id": 135,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        578,
        947
      ],
      [
        830,
        1177
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/scalebar_widget",
    "scrollable": false,
    "selected": false,
    "size": "252*230",
    "temp_id": 136,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        861,
        989
      ],
      [
        1080,
        1219
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      138
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/on_map_action_button",
    "scrollable": false,
    "selected": false,
    "size": "219*230",
    "temp_id": 137,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        861,
        989
      ],
      [
        1080,
        1219
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      139
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 137,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "219*230",
    "temp_id": 138,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        892,
        1020
      ],
      [
        1039,
        1167
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageButton",
    "clickable": true,
    "content_description": "Directions",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 138,
    "resource_id": "com.google.android.apps.maps:id/on_map_directions_button",
    "scrollable": false,
    "selected": false,
    "size": "147*147",
    "temp_id": 139,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1080,
        1000
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      141
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/on_map_secondary_action_button_container",
    "scrollable": false,
    "selected": false,
    "size": "199*199",
    "temp_id": 140,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1080,
        987
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      142
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 140,
    "resource_id": "com.google.android.apps.maps:id/qu_mylocation_container",
    "scrollable": false,
    "selected": false,
    "size": "199*186",
    "temp_id": 141,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1080,
        987
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      143
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Location services disabled. Enable location services to re-center map to your location.",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 141,
    "resource_id": "com.google.android.apps.maps:id/mylocation_button",
    "scrollable": false,
    "selected": false,
    "size": "199*186",
    "temp_id": 142,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1049,
        969
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      144,
      146
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 142,
    "resource_id": "com.google.android.apps.maps:id/fab_icon",
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 143,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1049,
        969
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      145
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 143,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 144,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1049,
        969
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 144,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 145,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1049,
        969
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      147
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 143,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 146,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        801
      ],
      [
        1049,
        969
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 146,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 147,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 148,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 149,
    "text": null,
    "visible": false
  }
]
