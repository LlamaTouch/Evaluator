[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      1
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 1,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 2,
    "resource_id": "com.google.android.apps.nexuslauncher:id/launcher",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      5,
      6,
      23,
      24,
      25
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 3,
    "resource_id": "com.google.android.apps.nexuslauncher:id/drag_layer",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/scrim_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      7,
      17
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/workspace",
    "scrollable": true,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        63
      ],
      [
        1030,
        1409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 6,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "980*1346",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        63
      ],
      [
        1030,
        1409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      9,
      16
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 7,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "980*1346",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        63
      ],
      [
        1030,
        303
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 8,
    "resource_id": "com.google.android.apps.nexuslauncher:id/search_container_workspace",
    "scrollable": false,
    "selected": false,
    "size": "980*240",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        64
      ],
      [
        1030,
        303
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 9,
    "resource_id": "com.google.android.apps.nexuslauncher:id/bc_smartspace_view",
    "scrollable": false,
    "selected": false,
    "size": "938*239",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        64
      ],
      [
        1030,
        303
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      12
    ],
    "class": "androidx.viewpager.widget.ViewPager",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 10,
    "resource_id": "com.google.android.apps.nexuslauncher:id/smartspace_card_pager",
    "scrollable": false,
    "selected": false,
    "size": "938*239",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        64
      ],
      [
        1030,
        303
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      13
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 11,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "938*239",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        100
      ],
      [
        1030,
        216
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      14,
      15
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 12,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "938*116",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        100
      ],
      [
        1030,
        155
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "Sun, Jan 21",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 13,
    "resource_id": "com.google.android.apps.nexuslauncher:id/clock",
    "scrollable": false,
    "selected": false,
    "size": "938*55",
    "temp_id": 14,
    "text": "Sun, Jan 21",
    "visible": true
  },
  {
    "bounds": [
      [
        92,
        173
      ],
      [
        92,
        216
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 13,
    "resource_id": "com.google.android.apps.nexuslauncher:id/subtitle_text",
    "scrollable": false,
    "selected": false,
    "size": "0*43",
    "temp_id": 15,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        50,
        615
      ],
      [
        268,
        855
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Maps",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "218*240",
    "temp_id": 16,
    "text": "Maps",
    "visible": true
  },
  {
    "bounds": [
      [
        1081,
        63
      ],
      [
        1080,
        1409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 6,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-1*1346",
    "temp_id": 17,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1081,
        63
      ],
      [
        1080,
        1409
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      19,
      20,
      21,
      22
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-1*1346",
    "temp_id": 18,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1589,
        891
      ],
      [
        1080,
        1131
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Play Store",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-509*240",
    "temp_id": 19,
    "text": "Play Store",
    "visible": false
  },
  {
    "bounds": [
      [
        1843,
        891
      ],
      [
        1080,
        1131
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Photos",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-763*240",
    "temp_id": 20,
    "text": "Photos",
    "visible": false
  },
  {
    "bounds": [
      [
        1589,
        1167
      ],
      [
        1080,
        1407
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Gmail",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-509*240",
    "temp_id": 21,
    "text": "Gmail",
    "visible": false
  },
  {
    "bounds": [
      [
        1843,
        1167
      ],
      [
        1080,
        1407
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "YouTube",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-763*240",
    "temp_id": 22,
    "text": "YouTube",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Home",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1729",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1377
      ],
      [
        1080,
        1440
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/page_indicator",
    "scrollable": false,
    "selected": false,
    "size": "1080*63",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1440
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      26,
      29
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/hotseat",
    "scrollable": false,
    "selected": false,
    "size": "1080*478",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        51,
        1440
      ],
      [
        1029,
        1609
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      27,
      28
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "978*169",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        306,
        1440
      ],
      [
        520,
        1609
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Messages",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "214*169",
    "temp_id": 27,
    "text": "Messages",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1440
      ],
      [
        775,
        1609
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Chrome",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "214*169",
    "temp_id": 28,
    "text": "Chrome",
    "visible": true
  },
  {
    "bounds": [
      [
        90,
        1622
      ],
      [
        990,
        1787
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      30,
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Search",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "900*165",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        132,
        1673
      ],
      [
        195,
        1736
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 29,
    "resource_id": "com.google.android.apps.nexuslauncher:id/g_icon",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        848,
        1622
      ],
      [
        990,
        1787
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 29,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "142*165",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        848,
        1622
      ],
      [
        990,
        1787
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 31,
    "resource_id": "com.google.android.apps.nexuslauncher:id/mic_icon",
    "scrollable": false,
    "selected": false,
    "size": "142*165",
    "temp_id": 32,
    "text": null,
    "visible": true
  }
]
