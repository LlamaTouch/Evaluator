[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      1
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 1,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 2,
    "resource_id": "com.google.android.apps.nexuslauncher:id/launcher",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      5,
      6,
      35,
      36,
      37
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 3,
    "resource_id": "com.google.android.apps.nexuslauncher:id/drag_layer",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/scrim_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      7,
      17
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/workspace",
    "scrollable": true,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        165
      ],
      [
        -1,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 6,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-1*1524",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        165
      ],
      [
        -3,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      9,
      16
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 7,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-3*1524",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        165
      ],
      [
        -3,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 8,
    "resource_id": "com.google.android.apps.nexuslauncher:id/search_container_workspace",
    "scrollable": false,
    "selected": false,
    "size": "-3*272",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        166
      ],
      [
        -3,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 9,
    "resource_id": "com.google.android.apps.nexuslauncher:id/bc_smartspace_view",
    "scrollable": false,
    "selected": false,
    "size": "-3*271",
    "temp_id": 10,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        166
      ],
      [
        -3,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      12
    ],
    "class": "androidx.viewpager.widget.ViewPager",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 10,
    "resource_id": "com.google.android.apps.nexuslauncher:id/smartspace_card_pager",
    "scrollable": false,
    "selected": false,
    "size": "-3*271",
    "temp_id": 11,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        166
      ],
      [
        -3,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      13
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 11,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-3*271",
    "temp_id": 12,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        207
      ],
      [
        -3,
        339
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      14,
      15
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 12,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-3*132",
    "temp_id": 13,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        207
      ],
      [
        -3,
        269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "Tue, Feb 6",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 13,
    "resource_id": "com.google.android.apps.nexuslauncher:id/clock",
    "scrollable": false,
    "selected": false,
    "size": "-3*62",
    "temp_id": 14,
    "text": "Tue, Feb 6",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        290
      ],
      [
        -923,
        339
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 13,
    "resource_id": "com.google.android.apps.nexuslauncher:id/subtitle_text",
    "scrollable": false,
    "selected": false,
    "size": "-923*49",
    "temp_id": 15,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        791
      ],
      [
        -755,
        1063
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Maps",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "-755*272",
    "temp_id": 16,
    "text": "Maps",
    "visible": false
  },
  {
    "bounds": [
      [
        57,
        165
      ],
      [
        1023,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 6,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "966*1524",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        165
      ],
      [
        1021,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 16,
    "children": [
      19,
      20,
      21,
      22,
      23,
      24,
      25,
      26,
      27,
      28,
      29,
      30,
      31,
      32,
      33,
      34
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "962*1524",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        165
      ],
      [
        269,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Spotify",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 19,
    "text": "Spotify",
    "visible": true
  },
  {
    "bounds": [
      [
        310,
        165
      ],
      [
        520,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Amazon Shopping",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 20,
    "text": "Amazon Shopping",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        165
      ],
      [
        771,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "X",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 21,
    "text": "X",
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        165
      ],
      [
        1021,
        437
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Wallet",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "209*272",
    "temp_id": 22,
    "text": "Wallet",
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        478
      ],
      [
        269,
        750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Expedia",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 23,
    "text": "Expedia",
    "visible": true
  },
  {
    "bounds": [
      [
        310,
        478
      ],
      [
        520,
        750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Calculator",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 24,
    "text": "Calculator",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        478
      ],
      [
        771,
        750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Duolingo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 25,
    "text": "Duolingo",
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        478
      ],
      [
        1021,
        750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Facebook",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "209*272",
    "temp_id": 26,
    "text": "Facebook",
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        791
      ],
      [
        269,
        1063
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Play Books",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 27,
    "text": "Play Books",
    "visible": true
  },
  {
    "bounds": [
      [
        310,
        791
      ],
      [
        520,
        1063
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Uber Eats",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 28,
    "text": "Uber Eats",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        791
      ],
      [
        771,
        1063
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Podcasts",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 29,
    "text": "Podcasts",
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        1104
      ],
      [
        269,
        1376
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "News",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 30,
    "text": "News",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1104
      ],
      [
        771,
        1376
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Play Store",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 31,
    "text": "Play Store",
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        1104
      ],
      [
        1021,
        1376
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Photos",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "209*272",
    "temp_id": 32,
    "text": "Photos",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1417
      ],
      [
        771,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Gmail",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*272",
    "temp_id": 33,
    "text": "Gmail",
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        1417
      ],
      [
        1021,
        1689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "YouTube",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "209*272",
    "temp_id": 34,
    "text": "YouTube",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Home",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1728
      ],
      [
        1080,
        1791
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/page_indicator",
    "scrollable": false,
    "selected": false,
    "size": "1080*63",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1791
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      38,
      41
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 4,
    "resource_id": "com.google.android.apps.nexuslauncher:id/hotseat",
    "scrollable": false,
    "selected": false,
    "size": "1080*609",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        59,
        1791
      ],
      [
        1021,
        1986
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      39,
      40
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "962*195",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        310,
        1791
      ],
      [
        520,
        1986
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Messages",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*195",
    "temp_id": 39,
    "text": "Messages",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1791
      ],
      [
        771,
        1986
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": "Chrome",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "210*195",
    "temp_id": 40,
    "text": "Chrome",
    "visible": true
  },
  {
    "bounds": [
      [
        82,
        2070
      ],
      [
        997,
        2235
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      43
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Search",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": true,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "915*165",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        124,
        2121
      ],
      [
        187,
        2184
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 41,
    "resource_id": "com.google.android.apps.nexuslauncher:id/g_icon",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        855,
        2070
      ],
      [
        997,
        2235
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "142*165",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        855,
        2070
      ],
      [
        997,
        2235
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.nexuslauncher",
    "parent": 43,
    "resource_id": "com.google.android.apps.nexuslauncher:id/mic_icon",
    "scrollable": false,
    "selected": false,
    "size": "142*165",
    "temp_id": 44,
    "text": null,
    "visible": true
  }
]
