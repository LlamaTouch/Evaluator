[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      1,
      67,
      68
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2274",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 2,
    "resource_id": "com.duolingo:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      6,
      7,
      8,
      66
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 4,
    "resource_id": "com.duolingo:id/sessionRoot",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": "com.duolingo:id/rampUpLessonQuitContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": "com.duolingo:id/loadingIndicator",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      9,
      10,
      11,
      17,
      18
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": "com.duolingo:id/challengeContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*2211",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        0,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        0,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/hideForKeyboardHelper",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 10,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        231
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      12,
      13,
      14
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/headerContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*168",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        105
      ],
      [
        126,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/quitButton",
    "scrollable": false,
    "selected": false,
    "size": "84*84",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        168,
        126
      ],
      [
        870,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/progress",
    "scrollable": false,
    "selected": false,
    "size": "702*42",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        105
      ],
      [
        1038,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      15,
      16
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": "You have 5 hearts left",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/heartsIndicator",
    "scrollable": false,
    "selected": false,
    "size": "126*84",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        115
      ],
      [
        989,
        178
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 14,
    "resource_id": "com.duolingo:id/heartIndicatorIcon",
    "scrollable": false,
    "selected": false,
    "size": "77*63",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        989,
        105
      ],
      [
        1038,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 14,
    "resource_id": "com.duolingo:id/heartNumber",
    "scrollable": false,
    "selected": false,
    "size": "49*84",
    "temp_id": 16,
    "text": "5",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        105
      ],
      [
        1080,
        231
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/headerPlaceholder",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        231
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/element_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*2043",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        231
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      20,
      59,
      60
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2043",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        231
      ],
      [
        1080,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      21
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 19,
    "resource_id": "com.duolingo:id/elementContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*1822",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        231
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      22,
      27,
      33
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 20,
    "resource_id": "com.duolingo:id/challenge_select",
    "scrollable": false,
    "selected": false,
    "size": "996*1822",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        231
      ],
      [
        1038,
        404
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      23,
      26
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 21,
    "resource_id": "com.duolingo:id/header",
    "scrollable": false,
    "selected": false,
    "size": "996*173",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        231
      ],
      [
        323,
        294
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      24,
      25
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 22,
    "resource_id": "com.duolingo:id/challengeIndicator",
    "scrollable": false,
    "selected": false,
    "size": "281*63",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        231
      ],
      [
        105,
        294
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 23,
    "resource_id": "com.duolingo:id/indicator",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        126,
        240
      ],
      [
        323,
        286
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 23,
    "resource_id": "com.duolingo:id/label",
    "scrollable": false,
    "selected": false,
    "size": "197*46",
    "temp_id": 25,
    "text": "NEW WORD",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        326
      ],
      [
        1038,
        404
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 22,
    "resource_id": "com.duolingo:id/challengeInstruction",
    "scrollable": false,
    "selected": false,
    "size": "996*78",
    "temp_id": 26,
    "text": "Select the correct image",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        446
      ],
      [
        1038,
        572
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      28,
      29,
      31,
      32
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 21,
    "resource_id": "com.duolingo:id/prompt",
    "scrollable": false,
    "selected": false,
    "size": "996*126",
    "temp_id": 27,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        446
      ],
      [
        42,
        446
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 28,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        446
      ],
      [
        168,
        572
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 27,
    "resource_id": "com.duolingo:id/nonCharacterSpeakerView",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        74,
        446
      ],
      [
        136,
        567
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 29,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "62*121",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        446
      ],
      [
        393,
        541
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 27,
    "resource_id": "com.duolingo:id/hintablePrompt",
    "scrollable": false,
    "selected": false,
    "size": "351*95",
    "temp_id": 31,
    "text": "la femme",
    "visible": true
  },
  {
    "bounds": [
      [
        232,
        447
      ],
      [
        351,
        572
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "119*125",
    "temp_id": 32,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        614
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      34
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 21,
    "resource_id": "com.duolingo:id/selection",
    "scrollable": false,
    "selected": false,
    "size": "996*1439",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        614
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      35,
      41,
      47,
      53
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*1439",
    "temp_id": 34,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        614
      ],
      [
        519,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      36,
      37
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/option1",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        614
      ],
      [
        519,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 35,
    "resource_id": "com.duolingo:id/buttonSparklesViewStub",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        614
      ],
      [
        519,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      38
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 35,
    "resource_id": "com.duolingo:id/delegate",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        654
      ],
      [
        477,
        1269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      39,
      40
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 37,
    "resource_id": "com.duolingo:id/content",
    "scrollable": false,
    "selected": false,
    "size": "393*615",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        654
      ],
      [
        477,
        1210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 38,
    "resource_id": "com.duolingo:id/svg",
    "scrollable": false,
    "selected": false,
    "size": "393*556",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        1210
      ],
      [
        477,
        1269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 38,
    "resource_id": "com.duolingo:id/imageText",
    "scrollable": false,
    "selected": false,
    "size": "393*59",
    "temp_id": 40,
    "text": "the boy",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        614
      ],
      [
        1038,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      43
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/option2",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        614
      ],
      [
        1038,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 41,
    "resource_id": "com.duolingo:id/buttonSparklesViewStub",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        614
      ],
      [
        1038,
        1313
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 41,
    "resource_id": "com.duolingo:id/delegate",
    "scrollable": false,
    "selected": false,
    "size": "477*699",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        654
      ],
      [
        996,
        1269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      45,
      46
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 43,
    "resource_id": "com.duolingo:id/content",
    "scrollable": false,
    "selected": false,
    "size": "393*615",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        654
      ],
      [
        996,
        1210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 44,
    "resource_id": "com.duolingo:id/svg",
    "scrollable": false,
    "selected": false,
    "size": "393*556",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        1210
      ],
      [
        996,
        1269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 44,
    "resource_id": "com.duolingo:id/imageText",
    "scrollable": false,
    "selected": false,
    "size": "393*59",
    "temp_id": 46,
    "text": "one",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1355
      ],
      [
        519,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      48,
      49
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/option3",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 47,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1355
      ],
      [
        519,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 47,
    "resource_id": "com.duolingo:id/buttonSparklesViewStub",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1355
      ],
      [
        519,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      50
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 47,
    "resource_id": "com.duolingo:id/delegate",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 49,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        1395
      ],
      [
        477,
        2009
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      51,
      52
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 49,
    "resource_id": "com.duolingo:id/content",
    "scrollable": false,
    "selected": false,
    "size": "393*614",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        1395
      ],
      [
        477,
        1950
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 50,
    "resource_id": "com.duolingo:id/svg",
    "scrollable": false,
    "selected": false,
    "size": "393*555",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        1950
      ],
      [
        477,
        2009
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 50,
    "resource_id": "com.duolingo:id/imageText",
    "scrollable": false,
    "selected": false,
    "size": "393*59",
    "temp_id": 52,
    "text": "the girl",
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1355
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      54,
      55
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/option4",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 53,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1355
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 53,
    "resource_id": "com.duolingo:id/buttonSparklesViewStub",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        561,
        1355
      ],
      [
        1038,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 53,
    "resource_id": "com.duolingo:id/delegate",
    "scrollable": false,
    "selected": false,
    "size": "477*698",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        1395
      ],
      [
        996,
        2009
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      57,
      58
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 55,
    "resource_id": "com.duolingo:id/content",
    "scrollable": false,
    "selected": false,
    "size": "393*614",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        1395
      ],
      [
        996,
        1950
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 56,
    "resource_id": "com.duolingo:id/svg",
    "scrollable": false,
    "selected": false,
    "size": "393*555",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        603,
        1950
      ],
      [
        996,
        2009
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 56,
    "resource_id": "com.duolingo:id/imageText",
    "scrollable": false,
    "selected": false,
    "size": "393*59",
    "temp_id": 58,
    "text": "the woman",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        444
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 19,
    "resource_id": "com.duolingo:id/gradingRibbonContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*1830",
    "temp_id": 59,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2095
      ],
      [
        1080,
        2232
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      61
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 19,
    "resource_id": "com.duolingo:id/buttonsContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*137",
    "temp_id": 60,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        2095
      ],
      [
        1038,
        2232
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      62,
      64
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 60,
    "resource_id": "com.duolingo:id/buttonsContainer",
    "scrollable": false,
    "selected": false,
    "size": "996*137",
    "temp_id": 61,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        2095
      ],
      [
        1038,
        2095
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      63
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*0",
    "temp_id": 62,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2095
      ],
      [
        1038,
        2095
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 62,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*0",
    "temp_id": 63,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2095
      ],
      [
        1038,
        2232
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      65
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 61,
    "resource_id": "com.duolingo:id/submitAndSkipContainer",
    "scrollable": false,
    "selected": false,
    "size": "996*137",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        2095
      ],
      [
        1038,
        2232
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": false,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 64,
    "resource_id": "com.duolingo:id/submitButton",
    "scrollable": false,
    "selected": false,
    "size": "996*137",
    "temp_id": 65,
    "text": "CHECK",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1099
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1175",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 0,
    "resource_id": "android:id/statusBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*63",
    "temp_id": 67,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2274
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 68,
    "text": null,
    "visible": false
  }
]
