[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      104
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      6
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      7
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      8,
      9,
      13
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/og_dialog_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 7,
    "resource_id": "com.google.android.apps.maps:id/og_dialog_scrim_ve",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      10,
      11
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 7,
    "resource_id": "com.google.android.apps.maps:id/og_container_header",
    "scrollable": false,
    "selected": false,
    "size": "1080*147",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        147,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Close",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 9,
    "resource_id": "com.google.android.apps.maps:id/og_header_close_button",
    "scrollable": false,
    "selected": false,
    "size": "147*147",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        147,
        105
      ],
      [
        933,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      12
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 9,
    "resource_id": "com.google.android.apps.maps:id/og_header_container",
    "scrollable": false,
    "selected": false,
    "size": "786*63",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        147,
        105
      ],
      [
        933,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 11,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "786*63",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 7,
    "resource_id": "com.google.android.apps.maps:id/og_container_scroll_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*1582",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1582",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      16,
      98,
      99
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": "com.google.android.apps.maps:id/og_container_scroll_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1582",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1080,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      17
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": "com.google.android.apps.maps:id/og_container_content_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1540",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1080,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      18,
      76
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": "com.google.android.apps.maps:id/og_has_selected_content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1540",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        210
      ],
      [
        1017,
        1354
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "androidx.cardview.widget.CardView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "954*1144",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        210
      ],
      [
        1017,
        1354
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      20,
      30,
      32,
      33
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "954*1144",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        210
      ],
      [
        1017,
        389
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      21,
      26,
      27,
      28
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/selected_account_view",
    "scrollable": false,
    "selected": false,
    "size": "954*179",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        231
      ],
      [
        231,
        368
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": "com.google.android.apps.maps:id/account_avatar_container",
    "scrollable": false,
    "selected": false,
    "size": "147*137",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        84,
        231
      ],
      [
        231,
        368
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      23,
      24,
      25
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Change profile picture.",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/account_avatar",
    "scrollable": false,
    "selected": false,
    "size": "147*137",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        89,
        231
      ],
      [
        89,
        231
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/badge_wrapper",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 23,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        89,
        231
      ],
      [
        89,
        231
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/ring_wrapper",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 24,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        89,
        231
      ],
      [
        226,
        368
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/og_apd_internal_image_view",
    "scrollable": false,
    "selected": false,
    "size": "137*137",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        245
      ],
      [
        295,
        303
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "Signed in as Ian\nagentian03@gmail.com",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": "com.google.android.apps.maps:id/og_primary_account_information",
    "scrollable": false,
    "selected": false,
    "size": "53*58",
    "temp_id": 26,
    "text": "Ian",
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        306
      ],
      [
        591,
        355
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": "com.google.android.apps.maps:id/og_secondary_account_information",
    "scrollable": false,
    "selected": false,
    "size": "349*49",
    "temp_id": 27,
    "text": "agentian03@gmail.com",
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        268
      ],
      [
        975,
        331
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": "com.google.android.apps.maps:id/og_trailing_drawable_container",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        268
      ],
      [
        975,
        331
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": "Expand account list.",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": "com.google.android.apps.maps:id/og_collapsed_chevron",
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        389
      ],
      [
        1017,
        515
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "954*126",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        389
      ],
      [
        828,
        515
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": "com.google.android.apps.maps:id/my_account_chip",
    "scrollable": false,
    "selected": false,
    "size": "586*126",
    "temp_id": 31,
    "text": "Manage your Google Account",
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        515
      ],
      [
        1017,
        557
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/og_top_cards",
    "scrollable": false,
    "selected": false,
    "size": "954*42",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        557
      ],
      [
        1017,
        1354
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 6,
    "children": [
      34,
      41,
      48,
      55,
      62,
      69
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/cards_and_actions",
    "scrollable": false,
    "selected": false,
    "size": "954*797",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        63,
        562
      ],
      [
        1017,
        694
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      35,
      40
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 34,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        594
      ],
      [
        975,
        694
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      36
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 34,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        599
      ],
      [
        975,
        689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      37
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        599
      ],
      [
        975,
        689
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      38,
      39
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        602
      ],
      [
        184,
        655
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        599
      ],
      [
        975,
        657
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 39,
    "text": "Turn on Incognito mode",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        628
      ],
      [
        975,
        628
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 34,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 40,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        63,
        694
      ],
      [
        1017,
        826
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      47
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        726
      ],
      [
        975,
        826
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        731
      ],
      [
        975,
        821
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      44
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 43,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        731
      ],
      [
        975,
        821
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      45,
      46
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 43,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        734
      ],
      [
        184,
        787
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        731
      ],
      [
        975,
        789
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 46,
    "text": "Your profile",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        760
      ],
      [
        975,
        760
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 47,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        63,
        826
      ],
      [
        1017,
        958
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      49,
      54
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        858
      ],
      [
        975,
        958
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      50
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 48,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 49,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        863
      ],
      [
        975,
        953
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      51
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 49,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        863
      ],
      [
        975,
        953
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      52,
      53
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 50,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        866
      ],
      [
        184,
        919
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 52,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        863
      ],
      [
        975,
        921
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 53,
    "text": "Your Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        892
      ],
      [
        975,
        892
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 48,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 54,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        63,
        958
      ],
      [
        1017,
        1090
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      56,
      61
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        990
      ],
      [
        975,
        1090
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      57
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        995
      ],
      [
        975,
        1085
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      58
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 56,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        995
      ],
      [
        975,
        1085
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      59,
      60
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 57,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        998
      ],
      [
        184,
        1051
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 59,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        995
      ],
      [
        975,
        1053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 60,
    "text": "Location sharing",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1024
      ],
      [
        975,
        1024
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 61,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        63,
        1090
      ],
      [
        1017,
        1222
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      63,
      68
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1122
      ],
      [
        975,
        1222
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      64
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 63,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1127
      ],
      [
        975,
        1217
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      65
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 63,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1127
      ],
      [
        975,
        1217
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      66,
      67
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1130
      ],
      [
        184,
        1183
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        1127
      ],
      [
        975,
        1185
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 67,
    "text": "Offline maps",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1156
      ],
      [
        975,
        1156
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 68,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        63,
        1222
      ],
      [
        1017,
        1354
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      70,
      75
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "954*132",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1254
      ],
      [
        975,
        1354
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      71
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1259
      ],
      [
        975,
        1349
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      72
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 71,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1259
      ],
      [
        975,
        1349
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      73,
      74
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 71,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1262
      ],
      [
        184,
        1315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 72,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 73,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        1259
      ],
      [
        975,
        1317
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 72,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 74,
    "text": "Add your business",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1288
      ],
      [
        975,
        1288
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 75,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1354
      ],
      [
        1080,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      77,
      84,
      91
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": "com.google.android.apps.maps:id/common_actions",
    "scrollable": false,
    "selected": false,
    "size": "1080*396",
    "temp_id": 76,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1354
      ],
      [
        1080,
        1486
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      78,
      83
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 76,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "1080*132",
    "temp_id": 77,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1386
      ],
      [
        975,
        1486
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      79
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 78,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1391
      ],
      [
        975,
        1481
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      80
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 78,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 79,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1391
      ],
      [
        975,
        1481
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      81,
      82
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 79,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 80,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1394
      ],
      [
        184,
        1447
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 81,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        1391
      ],
      [
        975,
        1449
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 82,
    "text": "Your data in Maps",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1420
      ],
      [
        975,
        1420
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 83,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1486
      ],
      [
        1080,
        1618
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      85,
      90
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 76,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "1080*132",
    "temp_id": 84,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1518
      ],
      [
        975,
        1618
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      86
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 84,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 85,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1523
      ],
      [
        975,
        1613
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      87
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 85,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 86,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1523
      ],
      [
        975,
        1613
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      88,
      89
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 86,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 87,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1526
      ],
      [
        184,
        1579
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 87,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 88,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        1523
      ],
      [
        975,
        1581
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 87,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 89,
    "text": "Settings",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1552
      ],
      [
        975,
        1552
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 84,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 90,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1618
      ],
      [
        1080,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      92,
      97
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 76,
    "resource_id": "com.google.android.apps.maps:id/og_card",
    "scrollable": false,
    "selected": false,
    "size": "1080*132",
    "temp_id": 91,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1650
      ],
      [
        975,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      93
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 91,
    "resource_id": "com.google.android.apps.maps:id/og_card_content_root",
    "scrollable": false,
    "selected": false,
    "size": "844*100",
    "temp_id": 92,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1655
      ],
      [
        975,
        1745
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      94
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 92,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 93,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1655
      ],
      [
        975,
        1745
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      95,
      96
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 93,
    "resource_id": "com.google.android.apps.maps:id/og_full_text_card_root",
    "scrollable": false,
    "selected": false,
    "size": "844*90",
    "temp_id": 94,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        131,
        1658
      ],
      [
        184,
        1711
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 94,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_icon",
    "scrollable": false,
    "selected": false,
    "size": "53*53",
    "temp_id": 95,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        242,
        1655
      ],
      [
        975,
        1713
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 94,
    "resource_id": "com.google.android.apps.maps:id/og_text_card_title",
    "scrollable": false,
    "selected": false,
    "size": "733*58",
    "temp_id": 96,
    "text": "Help & feedback",
    "visible": true
  },
  {
    "bounds": [
      [
        975,
        1684
      ],
      [
        975,
        1684
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 91,
    "resource_id": "com.google.android.apps.maps:id/og_highlight_container",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 97,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1750
      ],
      [
        1080,
        1750
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 98,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        163,
        1750
      ],
      [
        917,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      100
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": "com.google.android.apps.maps:id/og_container_footer",
    "scrollable": false,
    "selected": false,
    "size": "754*42",
    "temp_id": 99,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        163,
        1750
      ],
      [
        917,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      101,
      102,
      103
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 99,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "754*42",
    "temp_id": 100,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        226,
        1750
      ],
      [
        492,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 100,
    "resource_id": "com.google.android.apps.maps:id/og_privacy_policy_button",
    "scrollable": false,
    "selected": false,
    "size": "266*42",
    "temp_id": 101,
    "text": "Privacy Policy",
    "visible": true
  },
  {
    "bounds": [
      [
        513,
        1809
      ],
      [
        521,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 100,
    "resource_id": "com.google.android.apps.maps:id/og_separator1",
    "scrollable": false,
    "selected": false,
    "size": "8*-17",
    "temp_id": 102,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        542,
        1750
      ],
      [
        854,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 100,
    "resource_id": "com.google.android.apps.maps:id/og_tos_button",
    "scrollable": false,
    "selected": false,
    "size": "312*42",
    "temp_id": 103,
    "text": "Terms of Service",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 104,
    "text": null,
    "visible": false
  }
]
