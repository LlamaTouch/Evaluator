[
  {
    "bounds": [
      [
        28,
        459
      ],
      [
        1052,
        1333
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      1
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1024*874",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        28,
        459
      ],
      [
        1052,
        1333
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1024*874",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        28,
        459
      ],
      [
        1052,
        1333
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1024*874",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        28,
        459
      ],
      [
        1052,
        1333
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1024*874",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        501
      ],
      [
        1010,
        1291
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      5,
      6,
      7,
      8
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "940*790",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        501
      ],
      [
        1010,
        564
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "940*63",
    "temp_id": 5,
    "text": "Delete all Timeline data from this device?",
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        564
      ],
      [
        1010,
        999
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "940*435",
    "temp_id": 6,
    "text": "Your visits and routes will be deleted from your Timeline on this device. You may still have Timeline data saved on other devices or in Timeline backups.\n\nTo manage your Location History, visit Activity controls.",
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        999
      ],
      [
        1010,
        1125
      ]
    ],
    "checkable": true,
    "checked": true,
    "child_count": 0,
    "children": [],
    "class": "android.widget.CheckBox",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "940*126",
    "temp_id": 7,
    "text": "I understand and want to delete.",
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        1125
      ],
      [
        1010,
        1291
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      9,
      10,
      11
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "940*166",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        70,
        1151
      ],
      [
        563,
        1151
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "493*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        563,
        1151
      ],
      [
        791,
        1291
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "228*140",
    "temp_id": 10,
    "text": "Cancel",
    "visible": true
  },
  {
    "bounds": [
      [
        791,
        1151
      ],
      [
        1010,
        1291
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 8,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "219*140",
    "temp_id": 11,
    "text": "Delete",
    "visible": true
  }
]
