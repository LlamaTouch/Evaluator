[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      89
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 2,
    "resource_id": "com.duolingo:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      7
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": "com.duolingo:id/launchContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      8
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 5,
    "resource_id": "com.duolingo:id/homeContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*2400",
    "temp_id": 7,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 6,
    "children": [
      9,
      10,
      11,
      29,
      30,
      75
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 7,
    "resource_id": "com.duolingo:id/root",
    "scrollable": false,
    "selected": false,
    "size": "1080*2274",
    "temp_id": 8,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/homeLoadingIndicator",
    "scrollable": false,
    "selected": false,
    "size": "1080*2274",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/toolbarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*189",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      12,
      15,
      22,
      25,
      26
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/toolbar",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        165,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      13,
      14
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "Learning 2131888976",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/menuLanguage",
    "scrollable": false,
    "selected": false,
    "size": "165*126",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        165,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 12,
    "resource_id": "com.duolingo:id/itemButton",
    "scrollable": false,
    "selected": false,
    "size": "165*126",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        50,
        123
      ],
      [
        116,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 12,
    "resource_id": "com.duolingo:id/selectionMotionContainer",
    "scrollable": false,
    "selected": false,
    "size": "66*66",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        271,
        63
      ],
      [
        435,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      16,
      20,
      21
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "1 day streak",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/menuStreak",
    "scrollable": false,
    "selected": false,
    "size": "164*126",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        292,
        71
      ],
      [
        344,
        181
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      17,
      18
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 15,
    "resource_id": "com.duolingo:id/itemIconWrapper",
    "scrollable": false,
    "selected": false,
    "size": "52*110",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        292,
        95
      ],
      [
        344,
        158
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 16,
    "resource_id": "com.duolingo:id/imageView",
    "scrollable": false,
    "selected": false,
    "size": "52*63",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        292,
        95
      ],
      [
        344,
        158
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 16,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "52*63",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        292,
        95
      ],
      [
        344,
        158
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 18,
    "resource_id": "com.duolingo:id/shineView",
    "scrollable": false,
    "selected": false,
    "size": "52*63",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        320,
        123
      ],
      [
        386,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 15,
    "resource_id": "com.duolingo:id/selectionMotionContainer",
    "scrollable": false,
    "selected": false,
    "size": "66*66",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        365,
        63
      ],
      [
        435,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 15,
    "resource_id": "com.duolingo:id/itemButton",
    "scrollable": false,
    "selected": false,
    "size": "70*126",
    "temp_id": 21,
    "text": "1",
    "visible": true
  },
  {
    "bounds": [
      [
        540,
        63
      ],
      [
        777,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      23,
      24
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/menuShopV2",
    "scrollable": false,
    "selected": false,
    "size": "237*126",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        540,
        63
      ],
      [
        777,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 22,
    "resource_id": "com.duolingo:id/itemButton",
    "scrollable": false,
    "selected": false,
    "size": "237*126",
    "temp_id": 23,
    "text": "505",
    "visible": true
  },
  {
    "bounds": [
      [
        626,
        123
      ],
      [
        692,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 22,
    "resource_id": "com.duolingo:id/selectionMotionContainer",
    "scrollable": false,
    "selected": false,
    "size": "66*66",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        540,
        63
      ],
      [
        540,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/menuTitle",
    "scrollable": false,
    "selected": false,
    "size": "0*126",
    "temp_id": 25,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        883,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      27,
      28
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "You have 5 hearts left",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 11,
    "resource_id": "com.duolingo:id/menuCurrency",
    "scrollable": false,
    "selected": false,
    "size": "197*126",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        883,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 26,
    "resource_id": "com.duolingo:id/itemButton",
    "scrollable": false,
    "selected": false,
    "size": "197*126",
    "temp_id": 27,
    "text": "5",
    "visible": true
  },
  {
    "bounds": [
      [
        949,
        123
      ],
      [
        1015,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 26,
    "resource_id": "com.duolingo:id/selectionMotionContainer",
    "scrollable": false,
    "selected": false,
    "size": "66*66",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/drawerBackdrop",
    "scrollable": false,
    "selected": false,
    "size": "1080*2085",
    "temp_id": 29,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/fragmentContainerLearn",
    "scrollable": false,
    "selected": false,
    "size": "1080*1859",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 30,
    "resource_id": "com.duolingo:id/pathContainer",
    "scrollable": false,
    "selected": false,
    "size": "1080*1859",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      33,
      39
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1859",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      34
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 32,
    "resource_id": "com.duolingo:id/sectionHeader",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      35,
      36,
      37,
      38
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 34,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        189
      ],
      [
        1080,
        315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/sectionHeaderBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        189
      ],
      [
        105,
        315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/sectionMenu",
    "scrollable": false,
    "selected": false,
    "size": "63*126",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        349,
        223
      ],
      [
        731,
        282
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/sectionTitle",
    "scrollable": false,
    "selected": false,
    "size": "382*59",
    "temp_id": 37,
    "text": "Section\u00a01:\u00a0Rookie",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        310
      ],
      [
        1080,
        315
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 34,
    "resource_id": "com.duolingo:id/sectionHeaderBorder",
    "scrollable": false,
    "selected": false,
    "size": "1080*5",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        315
      ],
      [
        1080,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      40,
      45,
      53,
      69,
      72
    ],
    "class": "androidx.recyclerview.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 32,
    "resource_id": "com.duolingo:id/path",
    "scrollable": true,
    "selected": false,
    "size": "1080*1733",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        315
      ],
      [
        1080,
        557
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      41,
      42,
      43,
      44
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*242",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        315
      ],
      [
        1080,
        557
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 40,
    "resource_id": "com.duolingo:id/pathItemBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*242",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        357
      ],
      [
        901,
        435
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 40,
    "resource_id": "com.duolingo:id/title",
    "scrollable": false,
    "selected": false,
    "size": "859*78",
    "temp_id": 42,
    "text": "Unit 1",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        456
      ],
      [
        859,
        515
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 40,
    "resource_id": "com.duolingo:id/subtitle",
    "scrollable": false,
    "selected": false,
    "size": "817*59",
    "temp_id": 43,
    "text": "Use basic phrases, greet people",
    "visible": true
  },
  {
    "bounds": [
      [
        901,
        368
      ],
      [
        1038,
        505
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 40,
    "resource_id": "com.duolingo:id/guidebook",
    "scrollable": false,
    "selected": false,
    "size": "137*137",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        599
      ],
      [
        1080,
        974
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      46,
      50,
      51
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*375",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        441,
        599
      ],
      [
        643,
        767
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      47
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 45,
    "resource_id": "com.duolingo:id/tooltip",
    "scrollable": false,
    "selected": false,
    "size": "202*168",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        441,
        610
      ],
      [
        643,
        767
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      48
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 46,
    "resource_id": "com.duolingo:id/tooltip",
    "scrollable": false,
    "selected": false,
    "size": "202*157",
    "temp_id": 47,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        441,
        610
      ],
      [
        643,
        747
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      49
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 47,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "202*137",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        473,
        652
      ],
      [
        611,
        705
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 48,
    "resource_id": "com.duolingo:id/popupText",
    "scrollable": false,
    "selected": false,
    "size": "138*53",
    "temp_id": 49,
    "text": "START",
    "visible": true
  },
  {
    "bounds": [
      [
        412,
        730
      ],
      [
        669,
        974
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 45,
    "resource_id": "com.duolingo:id/progressRing",
    "scrollable": false,
    "selected": false,
    "size": "257*244",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        449,
        767
      ],
      [
        633,
        938
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      52
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 45,
    "resource_id": "com.duolingo:id/oval",
    "scrollable": false,
    "selected": false,
    "size": "184*171",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        449,
        767
      ],
      [
        633,
        928
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 51,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "184*161",
    "temp_id": 52,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        974
      ],
      [
        1080,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      54,
      63,
      65
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*781",
    "temp_id": 53,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        974
      ],
      [
        1080,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      55,
      58,
      61
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 53,
    "resource_id": "com.duolingo:id/item_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*781",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1030
      ],
      [
        1080,
        1201
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*171",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        331,
        1030
      ],
      [
        515,
        1201
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      57
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 55,
    "resource_id": "com.duolingo:id/oval",
    "scrollable": false,
    "selected": false,
    "size": "184*171",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        331,
        1030
      ],
      [
        515,
        1191
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 56,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "184*161",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1274
      ],
      [
        1080,
        1445
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      59
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*171",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        265,
        1274
      ],
      [
        449,
        1445
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      60
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 58,
    "resource_id": "com.duolingo:id/oval",
    "scrollable": false,
    "selected": false,
    "size": "184*171",
    "temp_id": 59,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        265,
        1274
      ],
      [
        449,
        1435
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 59,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "184*161",
    "temp_id": 60,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1519
      ],
      [
        1080,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      62
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*236",
    "temp_id": 61,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        318,
        1519
      ],
      [
        528,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 61,
    "resource_id": "com.duolingo:id/chest",
    "scrollable": false,
    "selected": false,
    "size": "210*236",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        527,
        974
      ],
      [
        1080,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      64
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 53,
    "resource_id": "com.duolingo:id/characterLottieAnimation",
    "scrollable": false,
    "selected": false,
    "size": "553*781",
    "temp_id": 63,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        527,
        974
      ],
      [
        1080,
        1755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 63,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "553*781",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        713,
        1528
      ],
      [
        894,
        1599
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      66,
      67,
      68
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 53,
    "resource_id": "com.duolingo:id/path_stars",
    "scrollable": false,
    "selected": false,
    "size": "181*71",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        713,
        1528
      ],
      [
        766,
        1578
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 65,
    "resource_id": "com.duolingo:id/star1",
    "scrollable": false,
    "selected": false,
    "size": "53*50",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        777,
        1549
      ],
      [
        830,
        1599
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 65,
    "resource_id": "com.duolingo:id/star2",
    "scrollable": false,
    "selected": false,
    "size": "53*50",
    "temp_id": 67,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        841,
        1528
      ],
      [
        894,
        1578
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 65,
    "resource_id": "com.duolingo:id/star3",
    "scrollable": false,
    "selected": false,
    "size": "53*50",
    "temp_id": 68,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1811
      ],
      [
        1080,
        1982
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      70
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*171",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        449,
        1811
      ],
      [
        633,
        1982
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      71
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 69,
    "resource_id": "com.duolingo:id/oval",
    "scrollable": false,
    "selected": false,
    "size": "184*171",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        449,
        1811
      ],
      [
        633,
        1972
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 70,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "184*161",
    "temp_id": 71,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2034
      ],
      [
        1080,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      73
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 39,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*14",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        567,
        2034
      ],
      [
        751,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      74
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 72,
    "resource_id": "com.duolingo:id/oval",
    "scrollable": false,
    "selected": false,
    "size": "184*14",
    "temp_id": 73,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        567,
        2034
      ],
      [
        751,
        2048
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 73,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "184*14",
    "temp_id": 74,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2048
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      76
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 8,
    "resource_id": "com.duolingo:id/tabs",
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 75,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2048
      ],
      [
        1080,
        2274
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 6,
    "children": [
      77,
      78,
      81,
      83,
      85,
      87
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 75,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*226",
    "temp_id": 76,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2048
      ],
      [
        1080,
        2053
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabBarBorder",
    "scrollable": false,
    "selected": false,
    "size": "1080*5",
    "temp_id": 77,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        75,
        2101
      ],
      [
        201,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      79,
      80
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "Learn Tab",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabLearn",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 78,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        75,
        2101
      ],
      [
        201,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 78,
    "resource_id": "com.duolingo:id/selectableBackground",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 79,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        88,
        2114
      ],
      [
        188,
        2214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 78,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "100*100",
    "temp_id": 80,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        276,
        2101
      ],
      [
        402,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      82
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "Leagues Tab",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabLeagues",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 81,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        289,
        2114
      ],
      [
        389,
        2214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 81,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "100*100",
    "temp_id": 82,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        477,
        2101
      ],
      [
        603,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      84
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "Profile Tab",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabProfile",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 83,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        490,
        2114
      ],
      [
        590,
        2214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 83,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "100*100",
    "temp_id": 84,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        678,
        2101
      ],
      [
        804,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      86
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "Goals Tab",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabGoals",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 85,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        691,
        2114
      ],
      [
        791,
        2214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 85,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "100*100",
    "temp_id": 86,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        879,
        2101
      ],
      [
        1005,
        2227
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      88
    ],
    "class": "android.view.ViewGroup",
    "clickable": true,
    "content_description": "News Tab",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 76,
    "resource_id": "com.duolingo:id/tabFeed",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 87,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        892,
        2114
      ],
      [
        992,
        2214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 87,
    "resource_id": "com.duolingo:id/icon",
    "scrollable": false,
    "selected": false,
    "size": "100*100",
    "temp_id": 88,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        2274
      ],
      [
        1080,
        2400
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.duolingo",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 89,
    "text": null,
    "visible": false
  }
]
