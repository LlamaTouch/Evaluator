[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      85
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      84
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 10,
    "children": [
      7,
      8,
      9,
      10,
      13,
      14,
      16,
      17,
      18,
      83
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        661
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      11
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1071*126",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        661
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      12
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 10,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1071*126",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        535
      ],
      [
        1071,
        535
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 11,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1071*0",
    "temp_id": 12,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 13,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/map_frame",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      20
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/fullscreen_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      21
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      23
    ],
    "class": "android.webkit.WebView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      24
    ],
    "class": "android.webkit.WebView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": true,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 23,
    "text": "Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      25
    ],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 23,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 24,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 24,
    "resource_id": "yDmH0d",
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 25,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      27
    ],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 25,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 26,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      28
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 27,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 28,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 29,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      31,
      53,
      63
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 29,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*1793",
    "temp_id": 30,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*336",
    "temp_id": 31,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      33,
      44
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*273",
    "temp_id": 32,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1084,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      34,
      35,
      37,
      40
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*147",
    "temp_id": 33,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        7,
        70
      ],
      [
        139,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 34,
    "text": "Back",
    "visible": true
  },
  {
    "bounds": [
      [
        126,
        105
      ],
      [
        958,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      36
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*63",
    "temp_id": 35,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        126,
        105
      ],
      [
        958,
        168
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*63",
    "temp_id": 36,
    "text": "Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        805,
        70
      ],
      [
        937,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      38
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 37,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        805,
        70
      ],
      [
        937,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      39
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 38,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        805,
        70
      ],
      [
        937,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*132",
    "temp_id": 39,
    "text": "Backup disabled.",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      41
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 40,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      42
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 41,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 42,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        945,
        70
      ],
      [
        1071,
        202
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*132",
    "temp_id": 43,
    "text": "More options",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      45
    ],
    "class": "android.widget.TabWidget",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*126",
    "temp_id": 44,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      46
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*126",
    "temp_id": 45,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        1084,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 6,
    "children": [
      47,
      48,
      49,
      50,
      51,
      52
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 45,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*126",
    "temp_id": 46,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        210
      ],
      [
        154,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab1",
    "scrollable": false,
    "selected": true,
    "size": "154*126",
    "temp_id": 47,
    "text": "Day",
    "visible": true
  },
  {
    "bounds": [
      [
        149,
        210
      ],
      [
        325,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab5",
    "scrollable": false,
    "selected": false,
    "size": "176*126",
    "temp_id": 48,
    "text": "Trips",
    "visible": true
  },
  {
    "bounds": [
      [
        320,
        210
      ],
      [
        546,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab6",
    "scrollable": false,
    "selected": false,
    "size": "226*126",
    "temp_id": 49,
    "text": "Insights",
    "visible": true
  },
  {
    "bounds": [
      [
        543,
        210
      ],
      [
        745,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab2",
    "scrollable": false,
    "selected": false,
    "size": "202*126",
    "temp_id": 50,
    "text": "Places",
    "visible": true
  },
  {
    "bounds": [
      [
        742,
        210
      ],
      [
        931,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab3",
    "scrollable": false,
    "selected": false,
    "size": "189*126",
    "temp_id": 51,
    "text": "Cities",
    "visible": true
  },
  {
    "bounds": [
      [
        926,
        210
      ],
      [
        1120,
        336
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": "tab4",
    "scrollable": false,
    "selected": false,
    "size": "194*126",
    "temp_id": 52,
    "text": "World",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        336
      ],
      [
        1084,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      54
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*561",
    "temp_id": 53,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        336
      ],
      [
        1084,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      55,
      59
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*561",
    "temp_id": 54,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        640,
        336
      ],
      [
        1084,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "444*160",
    "temp_id": 55,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        640,
        336
      ],
      [
        1084,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      57
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "444*160",
    "temp_id": 56,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        640,
        364
      ],
      [
        1042,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      58
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 56,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "402*132",
    "temp_id": 57,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        651,
        364
      ],
      [
        1029,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 57,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "378*132",
    "temp_id": 58,
    "text": "Timeline is on",
    "visible": true
  },
  {
    "bounds": [
      [
        868,
        748
      ],
      [
        1084,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      60
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "216*149",
    "temp_id": 59,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        868,
        748
      ],
      [
        1084,
        897
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      61
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 59,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "216*149",
    "temp_id": 60,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        910,
        748
      ],
      [
        1042,
        876
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      62
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 60,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*128",
    "temp_id": 61,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        910,
        748
      ],
      [
        1042,
        876
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*128",
    "temp_id": 62,
    "text": "Past visits layer is off",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        895
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      64
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*898",
    "temp_id": 63,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        895
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      65,
      80
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 63,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1084*898",
    "temp_id": 64,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -1084,
        895
      ],
      [
        2163,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      66,
      67,
      68
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "3247*898",
    "temp_id": 65,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -1063,
        947
      ],
      [
        -931,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "132*129",
    "temp_id": 66,
    "text": "Previous day",
    "visible": false
  },
  {
    "bounds": [
      [
        -149,
        947
      ],
      [
        -21,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "128*129",
    "temp_id": 67,
    "text": "Next day",
    "visible": false
  },
  {
    "bounds": [
      [
        -2,
        895
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      69,
      77
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*898",
    "temp_id": 68,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -2,
        895
      ],
      [
        1084,
        1097
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      70
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 68,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*202",
    "temp_id": 69,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -2,
        895
      ],
      [
        1084,
        1097
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      71,
      72,
      76
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*202",
    "temp_id": 70,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        506,
        916
      ],
      [
        574,
        929
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "68*13",
    "temp_id": 71,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -2,
        895
      ],
      [
        1084,
        1097
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      73,
      75
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*202",
    "temp_id": 72,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        18,
        947
      ],
      [
        147,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      74
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 72,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "129*129",
    "temp_id": 73,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        18,
        947
      ],
      [
        147,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 73,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "129*129",
    "temp_id": 74,
    "text": "Previous day",
    "visible": true
  },
  {
    "bounds": [
      [
        448,
        947
      ],
      [
        632,
        1076
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 72,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "184*129",
    "temp_id": 75,
    "text": "Today",
    "visible": true
  },
  {
    "bounds": [
      [
        -2,
        895
      ],
      [
        1084,
        1097
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*202",
    "temp_id": 76,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        -2,
        1094
      ],
      [
        1084,
        1793
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      78,
      79
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 68,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1086*699",
    "temp_id": 77,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        241,
        1097
      ],
      [
        861,
        1538
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Image",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "620*441",
    "temp_id": 78,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        349,
        1540
      ],
      [
        753,
        1596
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "404*56",
    "temp_id": 79,
    "text": "No visits for this day",
    "visible": true
  },
  {
    "bounds": [
      [
        897,
        1609
      ],
      [
        1050,
        1761
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      81
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "153*152",
    "temp_id": 80,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        897,
        1609
      ],
      [
        1050,
        1761
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      82
    ],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "153*152",
    "temp_id": 81,
    "text": "",
    "visible": true
  },
  {
    "bounds": [
      [
        897,
        1609
      ],
      [
        1050,
        1761
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 81,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "153*152",
    "temp_id": 82,
    "text": "Edit",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 83,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 84,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 85,
    "text": null,
    "visible": false
  }
]
