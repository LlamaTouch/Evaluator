[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      74
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      73
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 9,
    "children": [
      7,
      8,
      9,
      10,
      11,
      12,
      13,
      69,
      72
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 9,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 10,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      15
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": "com.google.android.apps.maps:id/fullscreen_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      16
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      17,
      27
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar",
    "scrollable": false,
    "selected": false,
    "size": "1080*211",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*148",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      20,
      21,
      24
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": "com.google.android.apps.maps:id/toolbar",
    "scrollable": false,
    "selected": false,
    "size": "1080*148",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1059,
        63
      ],
      [
        1059,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/end_section",
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 20,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        21,
        63
      ],
      [
        168,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/start_section",
    "scrollable": false,
    "selected": false,
    "size": "147*148",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        74
      ],
      [
        147,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      23
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Navigate up",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/nav_button",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        74
      ],
      [
        147,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar_button_icon",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        168,
        63
      ],
      [
        912,
        211
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      25
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": "com.google.android.apps.maps:id/title_frame",
    "scrollable": false,
    "selected": false,
    "size": "744*148",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        364,
        74
      ],
      [
        716,
        200
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      26
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 24,
    "resource_id": "com.google.android.apps.maps:id/title_section",
    "scrollable": false,
    "selected": false,
    "size": "352*126",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        364,
        103
      ],
      [
        716,
        171
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 25,
    "resource_id": "com.google.android.apps.maps:id/title",
    "scrollable": false,
    "selected": false,
    "size": "352*68",
    "temp_id": 26,
    "text": "Personal content",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      28
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 16,
    "resource_id": "com.google.android.apps.maps:id/mod_app_bar_fullscreen_content_view",
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 27,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 27,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      30
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 29,
    "resource_id": "android:id/list_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        211
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 9,
    "children": [
      32,
      35,
      41,
      47,
      50,
      54,
      57,
      61,
      65
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*1581",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        253
      ],
      [
        1080,
        346
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      33
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        253
      ],
      [
        1038,
        346
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      34
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        274
      ],
      [
        1038,
        325
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 33,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 34,
    "text": "Your Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        346
      ],
      [
        1080,
        538
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      36,
      39
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*192",
    "temp_id": 35,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        346
      ],
      [
        874,
        538
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      37,
      38
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*192",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        388
      ],
      [
        335,
        445
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "293*57",
    "temp_id": 37,
    "text": "Timeline emails",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        445
      ],
      [
        759,
        496
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "717*51",
    "temp_id": 38,
    "text": "Get highlights of your Timeline in your inbox",
    "visible": true
  },
  {
    "bounds": [
      [
        874,
        346
      ],
      [
        1038,
        538
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      40
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 35,
    "resource_id": "android:id/widget_frame",
    "scrollable": false,
    "selected": false,
    "size": "164*192",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        916,
        406
      ],
      [
        1038,
        477
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Switch",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 39,
    "resource_id": "com.google.android.apps.maps:id/switchWidget",
    "scrollable": false,
    "selected": false,
    "size": "122*71",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        538
      ],
      [
        1080,
        730
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      42,
      45
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*192",
    "temp_id": 41,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        538
      ],
      [
        874,
        730
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      43,
      44
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "832*192",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        580
      ],
      [
        319,
        637
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "277*57",
    "temp_id": 43,
    "text": "Google Photos",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        637
      ],
      [
        653,
        688
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "611*51",
    "temp_id": 44,
    "text": "Show your Google Photos in Timeline",
    "visible": true
  },
  {
    "bounds": [
      [
        874,
        538
      ],
      [
        1038,
        730
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      46
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 41,
    "resource_id": "android:id/widget_frame",
    "scrollable": false,
    "selected": false,
    "size": "164*192",
    "temp_id": 45,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        916,
        598
      ],
      [
        1038,
        669
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Switch",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 45,
    "resource_id": "com.google.android.apps.maps:id/switchWidget",
    "scrollable": false,
    "selected": false,
    "size": "122*71",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        772
      ],
      [
        1080,
        865
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      48
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 47,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        772
      ],
      [
        1038,
        865
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      49
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 47,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        793
      ],
      [
        1038,
        844
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 48,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 49,
    "text": "App history",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        865
      ],
      [
        1080,
        1100
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      51
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 50,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        865
      ],
      [
        1038,
        1100
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      52,
      53
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 50,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        907
      ],
      [
        507,
        964
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "465*57",
    "temp_id": 52,
    "text": "Web & App Activity is off\u00a0",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        964
      ],
      [
        1038,
        1058
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 51,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 53,
    "text": "Allow features to work properly like Timeline and search suggestions",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1142
      ],
      [
        1080,
        1235
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      55
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*93",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1142
      ],
      [
        1038,
        1235
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      56
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*93",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1163
      ],
      [
        1038,
        1214
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "996*51",
    "temp_id": 56,
    "text": "Location settings",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1235
      ],
      [
        1080,
        1470
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      58
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1235
      ],
      [
        1038,
        1470
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      59,
      60
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 57,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1277
      ],
      [
        304,
        1334
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "262*57",
    "temp_id": 59,
    "text": "Location is on",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1334
      ],
      [
        1038,
        1428
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 60,
    "text": "Let this app know your location for things like directions, navigation and search",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1470
      ],
      [
        1080,
        1705
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      62
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*235",
    "temp_id": 61,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1470
      ],
      [
        1038,
        1705
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      63,
      64
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*235",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1512
      ],
      [
        300,
        1569
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "258*57",
    "temp_id": 63,
    "text": "Timeline is on",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1569
      ],
      [
        1038,
        1663
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "996*94",
    "temp_id": 64,
    "text": "Rediscover the places you've been and the routes you've traveled",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1705
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      66
    ],
    "class": "android.widget.LinearLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*87",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1705
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      67,
      68
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*87",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1747
      ],
      [
        476,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 66,
    "resource_id": "android:id/title",
    "scrollable": false,
    "selected": false,
    "size": "434*45",
    "temp_id": 67,
    "text": "Delete all Timeline data",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1804
      ],
      [
        911,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 66,
    "resource_id": "android:id/summary",
    "scrollable": false,
    "selected": false,
    "size": "869*-12",
    "temp_id": 68,
    "text": "Permanently delete visits and routes from this device",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      70
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        189
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      71
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 69,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        63
      ],
      [
        1080,
        63
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 70,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 71,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 73,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 74,
    "text": null,
    "visible": false
  }
]
