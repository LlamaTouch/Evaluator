[
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      1,
      250
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": -1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1918",
    "temp_id": 0,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      2
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 1,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      3
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 1,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 2,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      4
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 2,
    "resource_id": "com.google.android.apps.maps:id/action_bar_root",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 3,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      5
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 3,
    "resource_id": "android:id/content",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 4,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      6,
      249
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 4,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 5,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 15,
    "children": [
      7,
      8,
      9,
      11,
      12,
      13,
      51,
      52,
      222,
      223,
      235,
      236,
      239,
      240,
      241
    ],
    "class": "android.view.ViewGroup",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/mainmap_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 6,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        0
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_header_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 7,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        0,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/expandingscrollview_container",
    "scrollable": true,
    "selected": false,
    "size": "0*1792",
    "temp_id": 8,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      10
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/map_frame",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 9,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 9,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 10,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/sidequest_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 11,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/fullscreens_group",
    "scrollable": false,
    "selected": false,
    "size": "1080*1792",
    "temp_id": 12,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      14
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*375",
    "temp_id": 13,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      15,
      36,
      50
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 13,
    "resource_id": "com.google.android.apps.maps:id/search_list_omnibox_layout",
    "scrollable": false,
    "selected": false,
    "size": "1080*375",
    "temp_id": 14,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        242
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      16,
      17
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*242",
    "temp_id": 15,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        242
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*242",
    "temp_id": 16,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        0
      ],
      [
        1080,
        242
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      18
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 15,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*242",
    "temp_id": 17,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        15,
        60
      ],
      [
        1065,
        234
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      19
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 17,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1050*174",
    "temp_id": 18,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      20
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 18,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 19,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      21
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 19,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 20,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      22
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 20,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 21,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      23,
      26,
      28,
      30,
      34
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 21,
    "resource_id": "com.google.android.apps.maps:id/mod_search_omnibox_layout",
    "scrollable": false,
    "selected": false,
    "size": "1018*126",
    "temp_id": 22,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        157,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      24
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 23,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        31,
        84
      ],
      [
        157,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      25
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Back",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 23,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_menu_button",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 24,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        62,
        115
      ],
      [
        125,
        178
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 24,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 25,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        84
      ],
      [
        797,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      27
    ],
    "class": "android.widget.EditText",
    "clickable": true,
    "content_description": "vegetarian restaurant",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_text_box",
    "scrollable": false,
    "selected": false,
    "size": "640*126",
    "temp_id": 26,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        157,
        84
      ],
      [
        797,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 26,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "640*126",
    "temp_id": 27,
    "text": "vegetarian restaurant",
    "visible": true
  },
  {
    "bounds": [
      [
        797,
        84
      ],
      [
        923,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      29
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_text_clear",
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 28,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        828,
        115
      ],
      [
        891,
        178
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": "Clear",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 28,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "63*63",
    "temp_id": 29,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        923,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      31
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 30,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        923,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      32
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 30,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 31,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        923,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      33
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 31,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 32,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        923,
        84
      ],
      [
        1049,
        210
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Voice search",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 32,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 33,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1049,
        147
      ],
      [
        1049,
        147
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      35
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 22,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 34,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1049,
        147
      ],
      [
        1049,
        147
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 34,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 35,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        221
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      37,
      48
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*154",
    "temp_id": 36,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        221
      ],
      [
        1080,
        367
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      38,
      40,
      42,
      44,
      46
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*146",
    "temp_id": 37,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        231
      ],
      [
        147,
        357
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      39
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "More filters",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 38,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        21,
        231
      ],
      [
        147,
        357
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "More filters",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 38,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 39,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        147,
        231
      ],
      [
        581,
        357
      ]
    ],
    "checkable": true,
    "checked": true,
    "child_count": 1,
    "children": [
      41
    ],
    "class": "android.widget.CompoundButton",
    "clickable": true,
    "content_description": "Vegetarian options",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "434*126",
    "temp_id": 40,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        147,
        231
      ],
      [
        581,
        357
      ]
    ],
    "checkable": true,
    "checked": true,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": false,
    "content_description": "Vegetarian options",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 40,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "434*126",
    "temp_id": 41,
    "text": "Vegetarian options",
    "visible": true
  },
  {
    "bounds": [
      [
        602,
        231
      ],
      [
        791,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 1,
    "children": [
      43
    ],
    "class": "android.widget.CompoundButton",
    "clickable": true,
    "content_description": "Dine-in",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "189*126",
    "temp_id": 42,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        602,
        231
      ],
      [
        791,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": false,
    "content_description": "Dine-in",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 42,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "189*126",
    "temp_id": 43,
    "text": "Dine-in",
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        231
      ],
      [
        1014,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 1,
    "children": [
      45
    ],
    "class": "android.widget.CompoundButton",
    "clickable": true,
    "content_description": "Takeout",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "202*126",
    "temp_id": 44,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        812,
        231
      ],
      [
        1014,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": false,
    "content_description": "Takeout",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 44,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "202*126",
    "temp_id": 45,
    "text": "Takeout",
    "visible": true
  },
  {
    "bounds": [
      [
        1035,
        231
      ],
      [
        1080,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 1,
    "children": [
      47
    ],
    "class": "android.widget.CompoundButton",
    "clickable": true,
    "content_description": "Delivery",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 37,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "45*126",
    "temp_id": 46,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1035,
        231
      ],
      [
        1080,
        357
      ]
    ],
    "checkable": true,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": false,
    "content_description": "Delivery",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 46,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "45*126",
    "temp_id": 47,
    "text": "Delivery",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      49
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 36,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*8",
    "temp_id": 48,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 48,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*8",
    "temp_id": 49,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 14,
    "resource_id": "com.google.android.apps.maps:id/search_omnibox_banner",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 50,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/home_bottom_sheet_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 51,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      53
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/custom_slider_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 52,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        367
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      54
    ],
    "class": "android.widget.ScrollView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 52,
    "resource_id": null,
    "scrollable": true,
    "selected": false,
    "size": "1080*1425",
    "temp_id": 53,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        723
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      55
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 53,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*1069",
    "temp_id": 54,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        723
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      56,
      58,
      139
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 54,
    "resource_id": "com.google.android.apps.maps:id/search_list_layout",
    "scrollable": true,
    "selected": false,
    "size": "1080*1069",
    "temp_id": 55,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        723
      ],
      [
        1080,
        755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      57
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*32",
    "temp_id": 56,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        723
      ],
      [
        1080,
        755
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 56,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*32",
    "temp_id": 57,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1647
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      59,
      83,
      84,
      120,
      123
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*892",
    "temp_id": 58,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      60
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*373",
    "temp_id": 59,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      61
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 59,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*373",
    "temp_id": 60,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      62
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 60,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*373",
    "temp_id": 61,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      63
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 61,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*373",
    "temp_id": 62,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        755
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      64
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 62,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*373",
    "temp_id": 63,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      65,
      71,
      77
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 63,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*352",
    "temp_id": 64,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        776
      ],
      [
        415,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      66
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 65,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        776
      ],
      [
        415,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      67
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 65,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 66,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        776
      ],
      [
        415,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      68
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 66,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 67,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        776
      ],
      [
        415,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      69,
      70
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 67,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 68,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        776
      ],
      [
        415,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 68,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 69,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        54,
        1090
      ],
      [
        78,
        1114
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 68,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "24*24",
    "temp_id": 70,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        776
      ],
      [
        809,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      72
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 71,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        776
      ],
      [
        809,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      73
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 71,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 72,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        776
      ],
      [
        809,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      74
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 72,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 73,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        776
      ],
      [
        809,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      75,
      76
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 73,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 74,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        776
      ],
      [
        809,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 74,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*352",
    "temp_id": 75,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        448,
        1090
      ],
      [
        472,
        1114
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 74,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "24*24",
    "temp_id": 76,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      78
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 64,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*352",
    "temp_id": 77,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      79
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 77,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*352",
    "temp_id": 78,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      80
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 78,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*352",
    "temp_id": 79,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      81,
      82
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 79,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*352",
    "temp_id": 80,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        776
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*352",
    "temp_id": 81,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        842,
        1090
      ],
      [
        866,
        1114
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 80,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "24*24",
    "temp_id": 82,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1080,
        1128
      ],
      [
        1080,
        1128
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 83,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1128
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      85,
      115
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*362",
    "temp_id": 84,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1159
      ],
      [
        1080,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      86,
      108
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 84,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*211",
    "temp_id": 85,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1159
      ],
      [
        912,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      87,
      89
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 85,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*211",
    "temp_id": 86,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1159
      ],
      [
        912,
        1217
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      88
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 86,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*58",
    "temp_id": 87,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1159
      ],
      [
        912,
        1217
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "Soul Vegetarian No. 2",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 87,
    "resource_id": "com.google.android.apps.maps:id/title",
    "scrollable": false,
    "selected": false,
    "size": "870*58",
    "temp_id": 88,
    "text": "Soul Vegetarian No. 2",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1217
      ],
      [
        912,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      90
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 86,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*153",
    "temp_id": 89,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1217
      ],
      [
        912,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      91,
      95,
      106
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 89,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*153",
    "temp_id": 90,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1217
      ],
      [
        418,
        1268
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      92
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 90,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*51",
    "temp_id": 91,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1217
      ],
      [
        418,
        1268
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      93,
      94
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 91,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*51",
    "temp_id": 92,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1217
      ],
      [
        418,
        1268
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 92,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*51",
    "temp_id": 93,
    "text": "4.3 stars (1,059)",
    "visible": true
  },
  {
    "bounds": [
      [
        418,
        1268
      ],
      [
        418,
        1268
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 92,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*0",
    "temp_id": 94,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        1268
      ],
      [
        912,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 7,
    "children": [
      96,
      97,
      98,
      101,
      102,
      104,
      105
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 90,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*51",
    "temp_id": 95,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1268
      ],
      [
        149,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "107*51",
    "temp_id": 96,
    "text": "Vegan",
    "visible": true
  },
  {
    "bounds": [
      [
        149,
        1268
      ],
      [
        179,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "30*51",
    "temp_id": 97,
    "text": " \u00b7 ",
    "visible": true
  },
  {
    "bounds": [
      [
        179,
        1268
      ],
      [
        313,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      99,
      100
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "134*51",
    "temp_id": 98,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        179,
        1268
      ],
      [
        180,
        1269
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 98,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1*1",
    "temp_id": 99,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        180,
        1268
      ],
      [
        313,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "$10 to $20",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 98,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "133*51",
    "temp_id": 100,
    "text": "$10\u201320",
    "visible": true
  },
  {
    "bounds": [
      [
        313,
        1268
      ],
      [
        343,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "30*51",
    "temp_id": 101,
    "text": " \u00b7 ",
    "visible": true
  },
  {
    "bounds": [
      [
        343,
        1268
      ],
      [
        912,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      103
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "569*51",
    "temp_id": 102,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        343,
        1268
      ],
      [
        912,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 102,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "569*51",
    "temp_id": 103,
    "text": "652 North Highland Avenue Northeast",
    "visible": true
  },
  {
    "bounds": [
      [
        907,
        1270
      ],
      [
        912,
        1317
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": "Wheelchair accessible",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "5*47",
    "temp_id": 104,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1268
      ],
      [
        912,
        1319
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 95,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*51",
    "temp_id": 105,
    "text": " \u00b7 ",
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        1319
      ],
      [
        518,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      107
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 90,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "476*51",
    "temp_id": 106,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1319
      ],
      [
        518,
        1370
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 106,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "476*51",
    "temp_id": 107,
    "text": "Closed \u00b7 Opens 1:00 PM\u00a0Tue",
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      109
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 85,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 108,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      110
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 108,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 109,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      111
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 109,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 110,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      112
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 110,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 111,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      113
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 111,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 112,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        912,
        1159
      ],
      [
        1038,
        1285
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      114
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Save Soul Vegetarian No. 2 to lists",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 112,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*126",
    "temp_id": 113,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        943,
        1164
      ],
      [
        1038,
        1259
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 113,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "95*95",
    "temp_id": 114,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1370
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      116
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 84,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*120",
    "temp_id": 115,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1370
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      117
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 115,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*120",
    "temp_id": 116,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1370
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      118
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 116,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*120",
    "temp_id": 117,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1385
      ],
      [
        1038,
        1483
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      119
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 117,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*98",
    "temp_id": 118,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        44,
        1387
      ],
      [
        1036,
        1481
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 118,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "992*94",
    "temp_id": 119,
    "text": "A Southern, meat-free menu (with gluten-free & vegan options) served in a casual space.",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1490
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      121
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 120,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1490
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      122
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 120,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 121,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1490
      ],
      [
        1080,
        1490
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 121,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 122,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1490
      ],
      [
        1080,
        1647
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      124
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 58,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 123,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1490
      ],
      [
        1080,
        1647
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      125
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 123,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 124,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1495
      ],
      [
        1038,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      126
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 124,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*126",
    "temp_id": 125,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1495
      ],
      [
        1038,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      127,
      130,
      133,
      136
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 125,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "996*126",
    "temp_id": 126,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1495
      ],
      [
        363,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      128
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 126,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*126",
    "temp_id": 127,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1495
      ],
      [
        363,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      129
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Directions to Soul Vegetarian No. 2, 652 North Highland Avenue Northeast",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 127,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*126",
    "temp_id": 128,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1505
      ],
      [
        363,
        1610
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Directions to Soul Vegetarian No. 2, 652 North Highland Avenue Northeast",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 128,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*105",
    "temp_id": 129,
    "text": "Directions",
    "visible": true
  },
  {
    "bounds": [
      [
        363,
        1495
      ],
      [
        745,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      131
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 126,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "382*126",
    "temp_id": 130,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        384,
        1495
      ],
      [
        745,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      132
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Order online",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 130,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "361*126",
    "temp_id": 131,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        384,
        1505
      ],
      [
        745,
        1610
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Order online",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 131,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "361*105",
    "temp_id": 132,
    "text": "Order online",
    "visible": true
  },
  {
    "bounds": [
      [
        745,
        1495
      ],
      [
        1006,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      134
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 126,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "261*126",
    "temp_id": 133,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        766,
        1495
      ],
      [
        1006,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      135
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Soul Vegetarian No. 2 Menu",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 133,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "240*126",
    "temp_id": 134,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        766,
        1505
      ],
      [
        1006,
        1610
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Soul Vegetarian No. 2 Menu",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 134,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "240*105",
    "temp_id": 135,
    "text": "Menu",
    "visible": true
  },
  {
    "bounds": [
      [
        1006,
        1495
      ],
      [
        1038,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      137
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 126,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "32*126",
    "temp_id": 136,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1027,
        1495
      ],
      [
        1038,
        1621
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      138
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Call Soul Vegetarian No. 2, 652 North Highland Avenue Northeast",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 136,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "11*126",
    "temp_id": 137,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        1027,
        1505
      ],
      [
        1038,
        1610
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Call Soul Vegetarian No. 2, 652 North Highland Avenue Northeast",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 137,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "11*105",
    "temp_id": 138,
    "text": "Call",
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 5,
    "children": [
      140,
      166,
      167,
      203,
      206
    ],
    "class": "android.widget.RelativeLayout",
    "clickable": true,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 55,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 139,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      141
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 139,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 140,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      142
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 140,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 141,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      143
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 141,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 142,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      144
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 142,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 143,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1668
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      145
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 143,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*124",
    "temp_id": 144,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      146,
      152,
      160
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 144,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "1080*103",
    "temp_id": 145,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1689
      ],
      [
        415,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      147
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 145,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 146,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1689
      ],
      [
        415,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      148
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 146,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 147,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1689
      ],
      [
        415,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      149
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 147,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 148,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1689
      ],
      [
        415,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      150,
      151
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 148,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 149,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        1689
      ],
      [
        415,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 149,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 150,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        54,
        2003
      ],
      [
        78,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 149,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "24*-211",
    "temp_id": 151,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      153
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 145,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 152,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      154
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 152,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 153,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      155
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 153,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 154,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      156
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Video",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 154,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 155,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      157
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 155,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 156,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      158,
      159
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 156,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 157,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 157,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 158,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        436,
        1689
      ],
      [
        809,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 157,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "373*103",
    "temp_id": 159,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      161
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 145,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*103",
    "temp_id": 160,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      162
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 160,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*103",
    "temp_id": 161,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      163
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 161,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*103",
    "temp_id": 162,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      164,
      165
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 162,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*103",
    "temp_id": 163,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        830,
        1689
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": true,
    "content_description": "Photo",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 163,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "250*103",
    "temp_id": 164,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        842,
        2003
      ],
      [
        866,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 163,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "24*-211",
    "temp_id": 165,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1080,
        2041
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 139,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*-249",
    "temp_id": 166,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2041
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      168,
      198
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 139,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-249",
    "temp_id": 167,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2072
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      169,
      191
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 167,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-280",
    "temp_id": 168,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2072
      ],
      [
        912,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      170,
      172
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 168,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*-280",
    "temp_id": 169,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2072
      ],
      [
        912,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      171
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 169,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*-280",
    "temp_id": 170,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2072
      ],
      [
        912,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "Green New American Vegetarian",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 170,
    "resource_id": "com.google.android.apps.maps:id/title",
    "scrollable": false,
    "selected": false,
    "size": "870*-280",
    "temp_id": 171,
    "text": "Green New American Vegetarian",
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2130
      ],
      [
        912,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      173
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 169,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*-338",
    "temp_id": 172,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2130
      ],
      [
        912,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 3,
    "children": [
      174,
      178,
      189
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 172,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "870*-338",
    "temp_id": 173,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2130
      ],
      [
        418,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      175
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 173,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*-338",
    "temp_id": 174,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2130
      ],
      [
        418,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      176,
      177
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 174,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*-338",
    "temp_id": 175,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2130
      ],
      [
        418,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 175,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "376*-338",
    "temp_id": 176,
    "text": "4.7 stars (2,520)",
    "visible": false
  },
  {
    "bounds": [
      [
        418,
        2181
      ],
      [
        418,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 175,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "0*-389",
    "temp_id": 177,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2181
      ],
      [
        641,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 7,
    "children": [
      179,
      180,
      181,
      184,
      185,
      187,
      188
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 173,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "599*-389",
    "temp_id": 178,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2181
      ],
      [
        149,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "107*-389",
    "temp_id": 179,
    "text": "Vegan",
    "visible": false
  },
  {
    "bounds": [
      [
        149,
        2181
      ],
      [
        179,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "30*-389",
    "temp_id": 180,
    "text": " \u00b7 ",
    "visible": false
  },
  {
    "bounds": [
      [
        179,
        2181
      ],
      [
        313,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      182,
      183
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "134*-389",
    "temp_id": 181,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        179,
        2181
      ],
      [
        180,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 181,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1*-389",
    "temp_id": 182,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        180,
        2181
      ],
      [
        313,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": "$10 to $20",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 181,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "133*-389",
    "temp_id": 183,
    "text": "$10\u201320",
    "visible": false
  },
  {
    "bounds": [
      [
        313,
        2181
      ],
      [
        343,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "30*-389",
    "temp_id": 184,
    "text": " \u00b7 ",
    "visible": false
  },
  {
    "bounds": [
      [
        343,
        2181
      ],
      [
        574,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      186
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*-389",
    "temp_id": 185,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        343,
        2181
      ],
      [
        574,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 185,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "231*-389",
    "temp_id": 186,
    "text": "2022 N 7th St",
    "visible": false
  },
  {
    "bounds": [
      [
        574,
        2181
      ],
      [
        604,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "30*-389",
    "temp_id": 187,
    "text": " \u00b7 ",
    "visible": false
  },
  {
    "bounds": [
      [
        599,
        2183
      ],
      [
        641,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": "Wheelchair accessible",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 178,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "42*-391",
    "temp_id": 188,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2232
      ],
      [
        469,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      190
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 173,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "427*-440",
    "temp_id": 189,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2232
      ],
      [
        469,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 189,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "427*-440",
    "temp_id": 190,
    "text": "Closed \u00b7 Opens 11:00 AM",
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      192
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 168,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 191,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      193
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 191,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 192,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      194
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 192,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 193,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      195
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 193,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 194,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      196
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 194,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 195,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        912,
        2072
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      197
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Save Green New American Vegetarian to lists",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 195,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "126*-280",
    "temp_id": 196,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        943,
        2077
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 196,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "95*-285",
    "temp_id": 197,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2283
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      199
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 167,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-491",
    "temp_id": 198,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2283
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      200
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 198,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-491",
    "temp_id": 199,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2283
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      201
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 199,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-491",
    "temp_id": 200,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2298
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      202
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 200,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*-506",
    "temp_id": 201,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        44,
        2300
      ],
      [
        1036,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.TextView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 201,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "992*-508",
    "temp_id": 202,
    "text": "Cheery restaurant turning out creative, vegan versions of familiar comfort foods.",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2403
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      204
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 139,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-611",
    "temp_id": 203,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2403
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      205
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 203,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-611",
    "temp_id": 204,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2403
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 204,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-611",
    "temp_id": 205,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2403
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      207
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 139,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-611",
    "temp_id": 206,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        2403
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      208
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 206,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*-611",
    "temp_id": 207,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2408
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      209
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 207,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "996*-616",
    "temp_id": 208,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2408
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 4,
    "children": [
      210,
      213,
      216,
      219
    ],
    "class": "android.support.v7.widget.RecyclerView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 208,
    "resource_id": "com.google.android.apps.maps:id/recycler_view",
    "scrollable": true,
    "selected": false,
    "size": "996*-616",
    "temp_id": 209,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2408
      ],
      [
        363,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      211
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 209,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*-616",
    "temp_id": 210,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2408
      ],
      [
        363,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      212
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Directions to Green New American Vegetarian, 2022 N 7th St",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 210,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*-616",
    "temp_id": 211,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        42,
        2418
      ],
      [
        363,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Directions to Green New American Vegetarian, 2022 N 7th St",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 211,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "321*-626",
    "temp_id": 212,
    "text": "Directions",
    "visible": false
  },
  {
    "bounds": [
      [
        363,
        2408
      ],
      [
        745,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      214
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 209,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "382*-616",
    "temp_id": 213,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        384,
        2408
      ],
      [
        745,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      215
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Order online",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 213,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "361*-616",
    "temp_id": 214,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        384,
        2418
      ],
      [
        745,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Order online",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 214,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "361*-626",
    "temp_id": 215,
    "text": "Order online",
    "visible": false
  },
  {
    "bounds": [
      [
        745,
        2408
      ],
      [
        1006,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      217
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 209,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "261*-616",
    "temp_id": 216,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        766,
        2408
      ],
      [
        1006,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      218
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Green New American Vegetarian Menu",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 216,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "240*-616",
    "temp_id": 217,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        766,
        2418
      ],
      [
        1006,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Green New American Vegetarian Menu",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 217,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "240*-626",
    "temp_id": 218,
    "text": "Menu",
    "visible": false
  },
  {
    "bounds": [
      [
        1006,
        2408
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      220
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 209,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "32*-616",
    "temp_id": 219,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1027,
        2408
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      221
    ],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Call Green New American Vegetarian, 2022 N 7th St",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 219,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "11*-616",
    "temp_id": 220,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        1027,
        2418
      ],
      [
        1038,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": "Call Green New American Vegetarian, 2022 N 7th St",
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 220,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "11*-626",
    "temp_id": 221,
    "text": "Call",
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        375
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/below_search_omnibox_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 222,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        663
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      224
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*288",
    "temp_id": 223,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        663
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      225
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 223,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*288",
    "temp_id": 224,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        532
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      226
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 224,
    "resource_id": "com.google.android.apps.maps:id/above_compass_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 225,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        375
      ],
      [
        1080,
        532
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      227
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 225,
    "resource_id": "com.google.android.apps.maps:id/layers_fab_button",
    "scrollable": false,
    "selected": false,
    "size": "1080*157",
    "temp_id": 226,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1080,
        532
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      228
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 226,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 227,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1080,
        532
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      229
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 227,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 228,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1080,
        532
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      230
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Layers",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 228,
    "resource_id": "com.google.android.apps.maps:id/layers_fab",
    "scrollable": false,
    "selected": false,
    "size": "152*142",
    "temp_id": 229,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1049,
        511
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      231,
      233
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 229,
    "resource_id": "com.google.android.apps.maps:id/fab_icon",
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 230,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1049,
        511
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      232
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 230,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 231,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1049,
        511
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 231,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 232,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1049,
        511
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      234
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 230,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 233,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        928,
        390
      ],
      [
        1049,
        511
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 233,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "121*121",
    "temp_id": 234,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        366,
        388
      ],
      [
        714,
        514
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/on_map_refresh_action_container",
    "scrollable": false,
    "selected": false,
    "size": "348*126",
    "temp_id": 235,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1562
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      237
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/footer_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*230",
    "temp_id": 236,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1562
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      238
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 236,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "1080*230",
    "temp_id": 237,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        669,
        1593
      ],
      [
        1039,
        1740
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.Button",
    "clickable": true,
    "content_description": "Map view",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 237,
    "resource_id": "com.google.android.apps.maps:id/map_list_toggle_fab",
    "scrollable": false,
    "selected": false,
    "size": "370*147",
    "temp_id": 238,
    "text": "View map",
    "visible": true
  },
  {
    "bounds": [
      [
        42,
        830
      ],
      [
        215,
        896
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/watermark_image",
    "scrollable": false,
    "selected": false,
    "size": "173*66",
    "temp_id": 239,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        598,
        681
      ],
      [
        850,
        880
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/scalebar_widget",
    "scrollable": false,
    "selected": false,
    "size": "252*199",
    "temp_id": 240,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1080,
        922
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      242
    ],
    "class": "android.widget.LinearLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 6,
    "resource_id": "com.google.android.apps.maps:id/on_map_secondary_action_button_container",
    "scrollable": false,
    "selected": false,
    "size": "199*199",
    "temp_id": 241,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1080,
        909
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      243
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 241,
    "resource_id": "com.google.android.apps.maps:id/qu_mylocation_container",
    "scrollable": false,
    "selected": false,
    "size": "199*186",
    "temp_id": 242,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1080,
        909
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      244
    ],
    "class": "android.widget.FrameLayout",
    "clickable": true,
    "content_description": "Location services disabled. Enable location services to re-center map to your location.",
    "editable": false,
    "enabled": true,
    "focusable": true,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 242,
    "resource_id": "com.google.android.apps.maps:id/mylocation_button",
    "scrollable": false,
    "selected": false,
    "size": "199*186",
    "temp_id": 243,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1049,
        891
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 2,
    "children": [
      245,
      247
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 243,
    "resource_id": "com.google.android.apps.maps:id/fab_icon",
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 244,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1049,
        891
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      246
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 244,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 245,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1049,
        891
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 245,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 246,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1049,
        891
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 1,
    "children": [
      248
    ],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 244,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 247,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        881,
        723
      ],
      [
        1049,
        891
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.ImageView",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 247,
    "resource_id": null,
    "scrollable": false,
    "selected": false,
    "size": "168*168",
    "temp_id": 248,
    "text": null,
    "visible": true
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1792
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.widget.FrameLayout",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 5,
    "resource_id": "com.google.android.apps.maps:id/survey_container",
    "scrollable": false,
    "selected": false,
    "size": "1080*0",
    "temp_id": 249,
    "text": null,
    "visible": false
  },
  {
    "bounds": [
      [
        0,
        1792
      ],
      [
        1080,
        1918
      ]
    ],
    "checkable": false,
    "checked": false,
    "child_count": 0,
    "children": [],
    "class": "android.view.View",
    "clickable": false,
    "content_description": null,
    "editable": false,
    "enabled": true,
    "focusable": false,
    "focused": false,
    "is_password": false,
    "long_clickable": false,
    "package": "com.google.android.apps.maps",
    "parent": 0,
    "resource_id": "android:id/navigationBarBackground",
    "scrollable": false,
    "selected": false,
    "size": "1080*126",
    "temp_id": 250,
    "text": null,
    "visible": false
  }
]
